module full_subber(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s,
  output       io_out_c
);
  wire [8:0] _result_T = io_in_a - io_in_b; // @[BinaryDesigns.scala 69:23]
  wire [9:0] _result_T_2 = _result_T - 9'h0; // @[BinaryDesigns.scala 69:34]
  wire [8:0] result = _result_T_2[8:0]; // @[BinaryDesigns.scala 68:22 69:12]
  assign io_out_s = result[7:0]; // @[BinaryDesigns.scala 70:23]
  assign io_out_c = result[8]; // @[BinaryDesigns.scala 71:23]
endmodule
module full_adder(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [23:0] io_out_s,
  output        io_out_c
);
  wire [24:0] _result_T = io_in_a + io_in_b; // @[BinaryDesigns.scala 55:23]
  wire [25:0] _result_T_1 = {{1'd0}, _result_T}; // @[BinaryDesigns.scala 55:34]
  wire [24:0] result = _result_T_1[24:0]; // @[BinaryDesigns.scala 54:22 55:12]
  assign io_out_s = result[23:0]; // @[BinaryDesigns.scala 56:23]
  assign io_out_c = result[24]; // @[BinaryDesigns.scala 57:23]
endmodule
module FP_adder_13ccs(
  input         clock,
  input         reset,
  input         io_in_en,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] subber_io_in_a; // @[FloatingPointDesigns.scala 1565:24]
  wire [7:0] subber_io_in_b; // @[FloatingPointDesigns.scala 1565:24]
  wire [7:0] subber_io_out_s; // @[FloatingPointDesigns.scala 1565:24]
  wire  subber_io_out_c; // @[FloatingPointDesigns.scala 1565:24]
  wire [23:0] adder_io_in_a; // @[FloatingPointDesigns.scala 1571:23]
  wire [23:0] adder_io_in_b; // @[FloatingPointDesigns.scala 1571:23]
  wire [23:0] adder_io_out_s; // @[FloatingPointDesigns.scala 1571:23]
  wire  adder_io_out_c; // @[FloatingPointDesigns.scala 1571:23]
  wire [7:0] subber2_io_in_a; // @[FloatingPointDesigns.scala 1632:25]
  wire [7:0] subber2_io_in_b; // @[FloatingPointDesigns.scala 1632:25]
  wire [7:0] subber2_io_out_s; // @[FloatingPointDesigns.scala 1632:25]
  wire  subber2_io_out_c; // @[FloatingPointDesigns.scala 1632:25]
  wire  sign_0 = io_in_a[31]; // @[FloatingPointDesigns.scala 1494:23]
  wire  sign_1 = io_in_b[31]; // @[FloatingPointDesigns.scala 1495:23]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FloatingPointDesigns.scala 1498:64]
  wire [8:0] _GEN_167 = {{1'd0}, io_in_a[30:23]}; // @[FloatingPointDesigns.scala 1498:36]
  wire [7:0] _GEN_0 = io_in_a[30:23] < 8'h1 ? 8'h1 : io_in_a[30:23]; // @[FloatingPointDesigns.scala 1500:46 1501:14 1503:14]
  wire [8:0] _GEN_1 = _GEN_167 > _T_2 ? _T_2 : {{1'd0}, _GEN_0}; // @[FloatingPointDesigns.scala 1498:71 1499:14]
  wire [8:0] _GEN_168 = {{1'd0}, io_in_b[30:23]}; // @[FloatingPointDesigns.scala 1505:36]
  wire [7:0] _GEN_2 = io_in_b[30:23] < 8'h1 ? 8'h1 : io_in_b[30:23]; // @[FloatingPointDesigns.scala 1507:45 1508:14 1510:14]
  wire [8:0] _GEN_3 = _GEN_168 > _T_2 ? _T_2 : {{1'd0}, _GEN_2}; // @[FloatingPointDesigns.scala 1505:71 1506:14]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FloatingPointDesigns.scala 1515:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FloatingPointDesigns.scala 1516:23]
  wire [23:0] whole_frac_0 = {1'h1,frac_0}; // @[FloatingPointDesigns.scala 1520:26]
  wire [23:0] whole_frac_1 = {1'h1,frac_1}; // @[FloatingPointDesigns.scala 1521:26]
  reg  sign_reg_0_0; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_0_1; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_1_0; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_1_1; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_2_0; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_2_1; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_3_0; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_3_1; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_4_0; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_4_1; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_5_0; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_5_1; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_6_0; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_6_1; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_7_0; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_7_1; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_8_0; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_8_1; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_9_0; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_9_1; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_10_0; // @[FloatingPointDesigns.scala 1523:28]
  reg  sign_reg_10_1; // @[FloatingPointDesigns.scala 1523:28]
  reg [7:0] exp_reg_0_0; // @[FloatingPointDesigns.scala 1524:28]
  reg [7:0] exp_reg_0_1; // @[FloatingPointDesigns.scala 1524:28]
  reg [7:0] exp_reg_1_0; // @[FloatingPointDesigns.scala 1524:28]
  reg [7:0] exp_reg_1_1; // @[FloatingPointDesigns.scala 1524:28]
  reg [7:0] exp_reg_2_0; // @[FloatingPointDesigns.scala 1524:28]
  reg [7:0] exp_reg_2_1; // @[FloatingPointDesigns.scala 1524:28]
  reg [22:0] frac_reg_0_0; // @[FloatingPointDesigns.scala 1525:28]
  reg [22:0] frac_reg_0_1; // @[FloatingPointDesigns.scala 1525:28]
  reg [22:0] frac_reg_1_0; // @[FloatingPointDesigns.scala 1525:28]
  reg [22:0] frac_reg_1_1; // @[FloatingPointDesigns.scala 1525:28]
  reg [22:0] frac_reg_2_0; // @[FloatingPointDesigns.scala 1525:28]
  reg [22:0] frac_reg_2_1; // @[FloatingPointDesigns.scala 1525:28]
  reg [23:0] wfrac_reg_0_0; // @[FloatingPointDesigns.scala 1526:28]
  reg [23:0] wfrac_reg_0_1; // @[FloatingPointDesigns.scala 1526:28]
  reg [23:0] wfrac_reg_1_0; // @[FloatingPointDesigns.scala 1526:28]
  reg [23:0] wfrac_reg_1_1; // @[FloatingPointDesigns.scala 1526:28]
  reg [23:0] wfrac_reg_2_0; // @[FloatingPointDesigns.scala 1526:28]
  reg [23:0] wfrac_reg_2_1; // @[FloatingPointDesigns.scala 1526:28]
  reg [7:0] subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1528:35]
  reg [7:0] subber_out_s_reg_1; // @[FloatingPointDesigns.scala 1528:35]
  reg  subber_out_c_reg_0; // @[FloatingPointDesigns.scala 1529:35]
  reg  subber_out_c_reg_1; // @[FloatingPointDesigns.scala 1529:35]
  reg [23:0] wire_temp_add_in_reg_0_0; // @[FloatingPointDesigns.scala 1531:39]
  reg [23:0] wire_temp_add_in_reg_0_1; // @[FloatingPointDesigns.scala 1531:39]
  reg [23:0] wire_temp_add_in_reg_1_0; // @[FloatingPointDesigns.scala 1531:39]
  reg [23:0] wire_temp_add_in_reg_1_1; // @[FloatingPointDesigns.scala 1531:39]
  reg  ref_s_reg_0; // @[FloatingPointDesigns.scala 1533:31]
  reg  ref_s_reg_1; // @[FloatingPointDesigns.scala 1533:31]
  reg  ref_s_reg_2; // @[FloatingPointDesigns.scala 1533:31]
  reg  ref_s_reg_3; // @[FloatingPointDesigns.scala 1533:31]
  reg  ref_s_reg_4; // @[FloatingPointDesigns.scala 1533:31]
  reg  ref_s_reg_5; // @[FloatingPointDesigns.scala 1533:31]
  reg  ref_s_reg_6; // @[FloatingPointDesigns.scala 1533:31]
  reg  ref_s_reg_7; // @[FloatingPointDesigns.scala 1533:31]
  reg [22:0] ref_frac_reg_0; // @[FloatingPointDesigns.scala 1534:31]
  reg [22:0] ref_frac_reg_1; // @[FloatingPointDesigns.scala 1534:31]
  reg [22:0] ref_frac_reg_2; // @[FloatingPointDesigns.scala 1534:31]
  reg [22:0] ref_frac_reg_3; // @[FloatingPointDesigns.scala 1534:31]
  reg [22:0] ref_frac_reg_4; // @[FloatingPointDesigns.scala 1534:31]
  reg [22:0] ref_frac_reg_5; // @[FloatingPointDesigns.scala 1534:31]
  reg [22:0] ref_frac_reg_6; // @[FloatingPointDesigns.scala 1534:31]
  reg [22:0] ref_frac_reg_7; // @[FloatingPointDesigns.scala 1534:31]
  reg [7:0] ref_exp_reg_0; // @[FloatingPointDesigns.scala 1535:31]
  reg [7:0] ref_exp_reg_1; // @[FloatingPointDesigns.scala 1535:31]
  reg [7:0] ref_exp_reg_2; // @[FloatingPointDesigns.scala 1535:31]
  reg [7:0] ref_exp_reg_3; // @[FloatingPointDesigns.scala 1535:31]
  reg [7:0] ref_exp_reg_4; // @[FloatingPointDesigns.scala 1535:31]
  reg [7:0] ref_exp_reg_5; // @[FloatingPointDesigns.scala 1535:31]
  reg [7:0] ref_exp_reg_6; // @[FloatingPointDesigns.scala 1535:31]
  reg [7:0] ref_exp_reg_7; // @[FloatingPointDesigns.scala 1535:31]
  reg [7:0] sub_exp_reg_0; // @[FloatingPointDesigns.scala 1536:31]
  reg [7:0] sub_exp_reg_1; // @[FloatingPointDesigns.scala 1536:31]
  reg [7:0] sub_exp_reg_2; // @[FloatingPointDesigns.scala 1536:31]
  reg [7:0] sub_exp_reg_3; // @[FloatingPointDesigns.scala 1536:31]
  reg [7:0] sub_exp_reg_4; // @[FloatingPointDesigns.scala 1536:31]
  reg [7:0] sub_exp_reg_5; // @[FloatingPointDesigns.scala 1536:31]
  reg [7:0] sub_exp_reg_6; // @[FloatingPointDesigns.scala 1536:31]
  reg [7:0] sub_exp_reg_7; // @[FloatingPointDesigns.scala 1536:31]
  reg [23:0] adder_io_out_s_reg_0; // @[FloatingPointDesigns.scala 1538:37]
  reg [23:0] adder_io_out_s_reg_1; // @[FloatingPointDesigns.scala 1538:37]
  reg [23:0] adder_io_out_s_reg_2; // @[FloatingPointDesigns.scala 1538:37]
  reg  adder_io_out_c_reg_0; // @[FloatingPointDesigns.scala 1539:37]
  reg  new_s_reg_0; // @[FloatingPointDesigns.scala 1541:35]
  reg  new_s_reg_1; // @[FloatingPointDesigns.scala 1541:35]
  reg  new_s_reg_2; // @[FloatingPointDesigns.scala 1541:35]
  reg  new_s_reg_3; // @[FloatingPointDesigns.scala 1541:35]
  reg  new_s_reg_4; // @[FloatingPointDesigns.scala 1541:35]
  reg  new_s_reg_5; // @[FloatingPointDesigns.scala 1541:35]
  reg [22:0] new_out_frac_reg_0; // @[FloatingPointDesigns.scala 1542:35]
  reg [7:0] new_out_exp_reg_0; // @[FloatingPointDesigns.scala 1543:35]
  reg  E_reg_0; // @[FloatingPointDesigns.scala 1544:24]
  reg  E_reg_1; // @[FloatingPointDesigns.scala 1544:24]
  reg  E_reg_2; // @[FloatingPointDesigns.scala 1544:24]
  reg  E_reg_3; // @[FloatingPointDesigns.scala 1544:24]
  reg  E_reg_4; // @[FloatingPointDesigns.scala 1544:24]
  reg  D_reg_0; // @[FloatingPointDesigns.scala 1545:24]
  reg  D_reg_1; // @[FloatingPointDesigns.scala 1545:24]
  reg  D_reg_2; // @[FloatingPointDesigns.scala 1545:24]
  reg  D_reg_3; // @[FloatingPointDesigns.scala 1545:24]
  reg  D_reg_4; // @[FloatingPointDesigns.scala 1545:24]
  reg [23:0] adder_result_reg_0; // @[FloatingPointDesigns.scala 1547:35]
  reg [23:0] adder_result_reg_1; // @[FloatingPointDesigns.scala 1547:35]
  reg [23:0] adder_result_reg_2; // @[FloatingPointDesigns.scala 1547:35]
  reg [5:0] leadingOne_reg_0; // @[FloatingPointDesigns.scala 1549:33]
  reg [5:0] leadingOne_reg_1; // @[FloatingPointDesigns.scala 1549:33]
  reg [31:0] io_in_a_reg_0; // @[FloatingPointDesigns.scala 1551:30]
  reg [31:0] io_in_a_reg_1; // @[FloatingPointDesigns.scala 1551:30]
  reg [31:0] io_in_a_reg_2; // @[FloatingPointDesigns.scala 1551:30]
  reg [31:0] io_in_a_reg_3; // @[FloatingPointDesigns.scala 1551:30]
  reg [31:0] io_in_a_reg_4; // @[FloatingPointDesigns.scala 1551:30]
  reg [31:0] io_in_a_reg_5; // @[FloatingPointDesigns.scala 1551:30]
  reg [31:0] io_in_a_reg_6; // @[FloatingPointDesigns.scala 1551:30]
  reg [31:0] io_in_a_reg_7; // @[FloatingPointDesigns.scala 1551:30]
  reg [31:0] io_in_a_reg_8; // @[FloatingPointDesigns.scala 1551:30]
  reg [31:0] io_in_a_reg_9; // @[FloatingPointDesigns.scala 1551:30]
  reg [31:0] io_in_a_reg_10; // @[FloatingPointDesigns.scala 1551:30]
  reg [31:0] io_in_b_reg_0; // @[FloatingPointDesigns.scala 1552:30]
  reg [31:0] io_in_b_reg_1; // @[FloatingPointDesigns.scala 1552:30]
  reg [31:0] io_in_b_reg_2; // @[FloatingPointDesigns.scala 1552:30]
  reg [31:0] io_in_b_reg_3; // @[FloatingPointDesigns.scala 1552:30]
  reg [31:0] io_in_b_reg_4; // @[FloatingPointDesigns.scala 1552:30]
  reg [31:0] io_in_b_reg_5; // @[FloatingPointDesigns.scala 1552:30]
  reg [31:0] io_in_b_reg_6; // @[FloatingPointDesigns.scala 1552:30]
  reg [31:0] io_in_b_reg_7; // @[FloatingPointDesigns.scala 1552:30]
  reg [31:0] io_in_b_reg_8; // @[FloatingPointDesigns.scala 1552:30]
  reg [31:0] io_in_b_reg_9; // @[FloatingPointDesigns.scala 1552:30]
  reg [31:0] io_in_b_reg_10; // @[FloatingPointDesigns.scala 1552:30]
  reg [7:0] subber2_out_s_reg_0; // @[FloatingPointDesigns.scala 1554:36]
  reg  subber2_out_c_reg_0; // @[FloatingPointDesigns.scala 1555:36]
  reg [7:0] cmpl_subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1576:40]
  wire [7:0] _cmpl_subber_out_s_reg_0_T = ~subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1578:41]
  wire [7:0] _cmpl_subber_out_s_reg_0_T_2 = 8'h1 + _cmpl_subber_out_s_reg_0_T; // @[FloatingPointDesigns.scala 1578:39]
  wire [23:0] _wire_temp_add_in_0_T = wfrac_reg_2_0 >> cmpl_subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1586:46]
  wire [23:0] _wire_temp_add_in_1_T = wfrac_reg_2_1 >> subber_out_s_reg_1; // @[FloatingPointDesigns.scala 1594:46]
  reg [23:0] cmpl_wire_temp_add_in_reg_0_0; // @[FloatingPointDesigns.scala 1597:44]
  reg [23:0] cmpl_wire_temp_add_in_reg_0_1; // @[FloatingPointDesigns.scala 1597:44]
  wire [23:0] _cmpl_wire_temp_add_in_reg_0_0_T = ~wire_temp_add_in_reg_0_0; // @[FloatingPointDesigns.scala 1599:48]
  wire [23:0] _cmpl_wire_temp_add_in_reg_0_0_T_2 = 24'h1 + _cmpl_wire_temp_add_in_reg_0_0_T; // @[FloatingPointDesigns.scala 1599:46]
  wire [23:0] _cmpl_wire_temp_add_in_reg_0_1_T = ~wire_temp_add_in_reg_0_1; // @[FloatingPointDesigns.scala 1600:48]
  wire [23:0] _cmpl_wire_temp_add_in_reg_0_1_T_2 = 24'h1 + _cmpl_wire_temp_add_in_reg_0_1_T; // @[FloatingPointDesigns.scala 1600:46]
  wire [1:0] _adder_io_in_a_T = {sign_reg_4_1,sign_reg_4_0}; // @[FloatingPointDesigns.scala 1603:38]
  wire  _new_s_T = ~adder_io_out_c_reg_0; // @[FloatingPointDesigns.scala 1610:15]
  wire  new_s = ~adder_io_out_c_reg_0 & (sign_reg_5_0 | sign_reg_5_1) | sign_reg_5_0 & sign_reg_5_1; // @[FloatingPointDesigns.scala 1610:75]
  wire  _D_T_1 = sign_reg_5_0 ^ sign_reg_5_1; // @[FloatingPointDesigns.scala 1617:53]
  wire  D = _new_s_T | sign_reg_5_0 ^ sign_reg_5_1; // @[FloatingPointDesigns.scala 1617:35]
  wire  E = _new_s_T & ~adder_io_out_s_reg_0[23] | _new_s_T & ~_D_T_1 | adder_io_out_c_reg_0 & adder_io_out_s_reg_0[23]
     & _D_T_1; // @[FloatingPointDesigns.scala 1619:134]
  reg [23:0] cmpl_adder_io_out_s_reg_0; // @[FloatingPointDesigns.scala 1621:42]
  wire [23:0] _cmpl_adder_io_out_s_reg_0_T = ~adder_io_out_s_reg_1; // @[FloatingPointDesigns.scala 1624:43]
  wire [23:0] _cmpl_adder_io_out_s_reg_0_T_2 = 24'h1 + _cmpl_adder_io_out_s_reg_0_T; // @[FloatingPointDesigns.scala 1624:41]
  wire [1:0] _adder_result_T = {sign_reg_7_1,sign_reg_7_0}; // @[FloatingPointDesigns.scala 1628:53]
  wire [1:0] _leadingOne_T_25 = adder_result_reg_0[2] ? 2'h2 : {{1'd0}, adder_result_reg_0[1]}; // @[FloatingPointDesigns.scala 1631:70]
  wire [1:0] _leadingOne_T_26 = adder_result_reg_0[3] ? 2'h3 : _leadingOne_T_25; // @[FloatingPointDesigns.scala 1631:70]
  wire [2:0] _leadingOne_T_27 = adder_result_reg_0[4] ? 3'h4 : {{1'd0}, _leadingOne_T_26}; // @[FloatingPointDesigns.scala 1631:70]
  wire [2:0] _leadingOne_T_28 = adder_result_reg_0[5] ? 3'h5 : _leadingOne_T_27; // @[FloatingPointDesigns.scala 1631:70]
  wire [2:0] _leadingOne_T_29 = adder_result_reg_0[6] ? 3'h6 : _leadingOne_T_28; // @[FloatingPointDesigns.scala 1631:70]
  wire [2:0] _leadingOne_T_30 = adder_result_reg_0[7] ? 3'h7 : _leadingOne_T_29; // @[FloatingPointDesigns.scala 1631:70]
  wire [3:0] _leadingOne_T_31 = adder_result_reg_0[8] ? 4'h8 : {{1'd0}, _leadingOne_T_30}; // @[FloatingPointDesigns.scala 1631:70]
  wire [3:0] _leadingOne_T_32 = adder_result_reg_0[9] ? 4'h9 : _leadingOne_T_31; // @[FloatingPointDesigns.scala 1631:70]
  wire [3:0] _leadingOne_T_33 = adder_result_reg_0[10] ? 4'ha : _leadingOne_T_32; // @[FloatingPointDesigns.scala 1631:70]
  wire [3:0] _leadingOne_T_34 = adder_result_reg_0[11] ? 4'hb : _leadingOne_T_33; // @[FloatingPointDesigns.scala 1631:70]
  wire [3:0] _leadingOne_T_35 = adder_result_reg_0[12] ? 4'hc : _leadingOne_T_34; // @[FloatingPointDesigns.scala 1631:70]
  wire [3:0] _leadingOne_T_36 = adder_result_reg_0[13] ? 4'hd : _leadingOne_T_35; // @[FloatingPointDesigns.scala 1631:70]
  wire [3:0] _leadingOne_T_37 = adder_result_reg_0[14] ? 4'he : _leadingOne_T_36; // @[FloatingPointDesigns.scala 1631:70]
  wire [3:0] _leadingOne_T_38 = adder_result_reg_0[15] ? 4'hf : _leadingOne_T_37; // @[FloatingPointDesigns.scala 1631:70]
  wire [4:0] _leadingOne_T_39 = adder_result_reg_0[16] ? 5'h10 : {{1'd0}, _leadingOne_T_38}; // @[FloatingPointDesigns.scala 1631:70]
  wire [4:0] _leadingOne_T_40 = adder_result_reg_0[17] ? 5'h11 : _leadingOne_T_39; // @[FloatingPointDesigns.scala 1631:70]
  wire [4:0] _leadingOne_T_41 = adder_result_reg_0[18] ? 5'h12 : _leadingOne_T_40; // @[FloatingPointDesigns.scala 1631:70]
  wire [4:0] _leadingOne_T_42 = adder_result_reg_0[19] ? 5'h13 : _leadingOne_T_41; // @[FloatingPointDesigns.scala 1631:70]
  wire [4:0] _leadingOne_T_43 = adder_result_reg_0[20] ? 5'h14 : _leadingOne_T_42; // @[FloatingPointDesigns.scala 1631:70]
  wire [4:0] _leadingOne_T_44 = adder_result_reg_0[21] ? 5'h15 : _leadingOne_T_43; // @[FloatingPointDesigns.scala 1631:70]
  wire [4:0] _leadingOne_T_45 = adder_result_reg_0[22] ? 5'h16 : _leadingOne_T_44; // @[FloatingPointDesigns.scala 1631:70]
  wire [4:0] _leadingOne_T_46 = adder_result_reg_0[23] ? 5'h17 : _leadingOne_T_45; // @[FloatingPointDesigns.scala 1631:70]
  wire [5:0] leadingOne = _leadingOne_T_46 + 5'h1; // @[FloatingPointDesigns.scala 1631:77]
  wire [5:0] _subber2_io_in_b_T_1 = 6'h18 - leadingOne_reg_0; // @[FloatingPointDesigns.scala 1634:42]
  wire [7:0] exp_0 = _GEN_1[7:0]; // @[FloatingPointDesigns.scala 1496:19]
  wire [7:0] exp_1 = _GEN_3[7:0]; // @[FloatingPointDesigns.scala 1496:19]
  reg [31:0] reg_out_s; // @[FloatingPointDesigns.scala 1705:28]
  wire [8:0] _GEN_169 = {{1'd0}, ref_exp_reg_7}; // @[FloatingPointDesigns.scala 1722:29]
  wire [23:0] _new_out_frac_reg_0_T_2 = 24'h800000 - 24'h1; // @[FloatingPointDesigns.scala 1724:60]
  wire [7:0] _new_out_exp_reg_0_T_3 = ref_exp_reg_7 + 8'h1; // @[FloatingPointDesigns.scala 1726:48]
  wire [8:0] _GEN_142 = _GEN_169 == _T_2 ? _T_2 : {{1'd0}, _new_out_exp_reg_0_T_3}; // @[FloatingPointDesigns.scala 1722:66 1723:30 1726:30]
  wire [23:0] _GEN_143 = _GEN_169 == _T_2 ? _new_out_frac_reg_0_T_2 : {{1'd0}, adder_result_reg_2[23:1]}; // @[FloatingPointDesigns.scala 1722:66 1724:31 1727:31]
  wire [5:0] _new_out_frac_reg_0_T_6 = 6'h18 - leadingOne_reg_1; // @[FloatingPointDesigns.scala 1740:94]
  wire [85:0] _GEN_5 = {{63'd0}, adder_result_reg_2[22:0]}; // @[FloatingPointDesigns.scala 1740:73]
  wire [85:0] _new_out_frac_reg_0_T_7 = _GEN_5 << _new_out_frac_reg_0_T_6; // @[FloatingPointDesigns.scala 1740:73]
  wire [7:0] _GEN_144 = subber2_out_c_reg_0 ? 8'h1 : subber2_out_s_reg_0; // @[FloatingPointDesigns.scala 1735:46 1736:32 1739:32]
  wire [85:0] _GEN_145 = subber2_out_c_reg_0 ? 86'h0 : _new_out_frac_reg_0_T_7; // @[FloatingPointDesigns.scala 1735:46 1737:33 1740:33]
  wire [7:0] _GEN_146 = leadingOne_reg_1 == 6'h1 & adder_result_reg_2 == 24'h0 & ((sign_reg_10_0 ^ sign_reg_10_1) &
    io_in_a_reg_10[30:0] == io_in_b_reg_10[30:0]) ? 8'h0 : _GEN_144; // @[FloatingPointDesigns.scala 1731:184 1732:30]
  wire [85:0] _GEN_147 = leadingOne_reg_1 == 6'h1 & adder_result_reg_2 == 24'h0 & ((sign_reg_10_0 ^ sign_reg_10_1) &
    io_in_a_reg_10[30:0] == io_in_b_reg_10[30:0]) ? 86'h0 : _GEN_145; // @[FloatingPointDesigns.scala 1731:184 1733:31]
  wire  _GEN_148 = D_reg_4 ? new_s_reg_4 : new_s_reg_5; // @[FloatingPointDesigns.scala 1729:36 1730:22 1541:35]
  wire [7:0] _GEN_149 = D_reg_4 ? _GEN_146 : new_out_exp_reg_0; // @[FloatingPointDesigns.scala 1543:35 1729:36]
  wire [85:0] _GEN_150 = D_reg_4 ? _GEN_147 : {{63'd0}, new_out_frac_reg_0}; // @[FloatingPointDesigns.scala 1542:35 1729:36]
  wire  _GEN_151 = ~D_reg_4 ? new_s_reg_4 : _GEN_148; // @[FloatingPointDesigns.scala 1720:36 1721:22]
  wire [8:0] _GEN_152 = ~D_reg_4 ? _GEN_142 : {{1'd0}, _GEN_149}; // @[FloatingPointDesigns.scala 1720:36]
  wire [85:0] _GEN_153 = ~D_reg_4 ? {{62'd0}, _GEN_143} : _GEN_150; // @[FloatingPointDesigns.scala 1720:36]
  wire  _GEN_154 = E_reg_4 ? new_s_reg_4 : _GEN_151; // @[FloatingPointDesigns.scala 1716:36 1717:22]
  wire [8:0] _GEN_155 = E_reg_4 ? {{1'd0}, ref_exp_reg_7} : _GEN_152; // @[FloatingPointDesigns.scala 1716:36 1718:28]
  wire [85:0] _GEN_156 = E_reg_4 ? {{63'd0}, adder_result_reg_2[22:0]} : _GEN_153; // @[FloatingPointDesigns.scala 1716:36 1719:29]
  wire [85:0] _GEN_158 = sub_exp_reg_7 >= 8'h17 ? {{63'd0}, ref_frac_reg_7} : _GEN_156; // @[FloatingPointDesigns.scala 1712:48 1714:29]
  wire [8:0] _GEN_159 = sub_exp_reg_7 >= 8'h17 ? {{1'd0}, ref_exp_reg_7} : _GEN_155; // @[FloatingPointDesigns.scala 1712:48 1715:28]
  wire [8:0] _GEN_161 = io_in_a_reg_10[30:0] == 31'h0 & io_in_b_reg_10[30:0] == 31'h0 ? 9'h0 : _GEN_159; // @[FloatingPointDesigns.scala 1708:86 1710:28]
  wire [85:0] _GEN_162 = io_in_a_reg_10[30:0] == 31'h0 & io_in_b_reg_10[30:0] == 31'h0 ? 86'h0 : _GEN_158; // @[FloatingPointDesigns.scala 1708:86 1711:29]
  wire [31:0] _reg_out_s_T_1 = {new_s_reg_5,new_out_exp_reg_0,new_out_frac_reg_0}; // @[FloatingPointDesigns.scala 1744:55]
  wire [8:0] _GEN_164 = io_in_en ? _GEN_161 : {{1'd0}, new_out_exp_reg_0}; // @[FloatingPointDesigns.scala 1707:20 1543:35]
  wire [85:0] _GEN_165 = io_in_en ? _GEN_162 : {{63'd0}, new_out_frac_reg_0}; // @[FloatingPointDesigns.scala 1707:20 1542:35]
  wire [85:0] _GEN_170 = reset ? 86'h0 : _GEN_165; // @[FloatingPointDesigns.scala 1542:{35,35}]
  wire [8:0] _GEN_171 = reset ? 9'h0 : _GEN_164; // @[FloatingPointDesigns.scala 1543:{35,35}]
  full_subber subber ( // @[FloatingPointDesigns.scala 1565:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  full_adder adder ( // @[FloatingPointDesigns.scala 1571:23]
    .io_in_a(adder_io_in_a),
    .io_in_b(adder_io_in_b),
    .io_out_s(adder_io_out_s),
    .io_out_c(adder_io_out_c)
  );
  full_subber subber2 ( // @[FloatingPointDesigns.scala 1632:25]
    .io_in_a(subber2_io_in_a),
    .io_in_b(subber2_io_in_b),
    .io_out_s(subber2_io_out_s),
    .io_out_c(subber2_io_out_c)
  );
  assign io_out_s = reg_out_s; // @[FloatingPointDesigns.scala 1706:14]
  assign subber_io_in_a = exp_reg_0_0; // @[FloatingPointDesigns.scala 1566:20]
  assign subber_io_in_b = exp_reg_0_1; // @[FloatingPointDesigns.scala 1567:20]
  assign adder_io_in_a = _adder_io_in_a_T == 2'h1 ? cmpl_wire_temp_add_in_reg_0_0 : wire_temp_add_in_reg_1_0; // @[FloatingPointDesigns.scala 1603:25]
  assign adder_io_in_b = _adder_io_in_a_T == 2'h2 ? cmpl_wire_temp_add_in_reg_0_1 : wire_temp_add_in_reg_1_1; // @[FloatingPointDesigns.scala 1604:25]
  assign subber2_io_in_a = ref_exp_reg_6; // @[FloatingPointDesigns.scala 1633:21]
  assign subber2_io_in_b = {{2'd0}, _subber2_io_in_b_T_1}; // @[FloatingPointDesigns.scala 1634:21]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_0_0 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_0_0 <= sign_0; // @[FloatingPointDesigns.scala 1642:19]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_0_1 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_0_1 <= sign_1; // @[FloatingPointDesigns.scala 1642:19]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_1_0 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_1_0 <= sign_reg_0_0; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_1_1 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_1_1 <= sign_reg_0_1; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_2_0 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_2_0 <= sign_reg_1_0; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_2_1 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_2_1 <= sign_reg_1_1; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_3_0 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_3_0 <= sign_reg_2_0; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_3_1 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_3_1 <= sign_reg_2_1; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_4_0 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_4_0 <= sign_reg_3_0; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_4_1 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_4_1 <= sign_reg_3_1; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_5_0 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_5_0 <= sign_reg_4_0; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_5_1 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_5_1 <= sign_reg_4_1; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_6_0 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_6_0 <= sign_reg_5_0; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_6_1 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_6_1 <= sign_reg_5_1; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_7_0 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_7_0 <= sign_reg_6_0; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_7_1 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_7_1 <= sign_reg_6_1; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_8_0 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_8_0 <= sign_reg_7_0; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_8_1 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_8_1 <= sign_reg_7_1; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_9_0 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_9_0 <= sign_reg_8_0; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_9_1 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_9_1 <= sign_reg_8_1; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_10_0 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_10_0 <= sign_reg_9_0; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1523:28]
      sign_reg_10_1 <= 1'h0; // @[FloatingPointDesigns.scala 1523:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sign_reg_10_1 <= sign_reg_9_1; // @[FloatingPointDesigns.scala 1675:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1524:28]
      exp_reg_0_0 <= 8'h0; // @[FloatingPointDesigns.scala 1524:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      exp_reg_0_0 <= exp_0; // @[FloatingPointDesigns.scala 1643:18]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1524:28]
      exp_reg_0_1 <= 8'h0; // @[FloatingPointDesigns.scala 1524:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      exp_reg_0_1 <= exp_1; // @[FloatingPointDesigns.scala 1643:18]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1524:28]
      exp_reg_1_0 <= 8'h0; // @[FloatingPointDesigns.scala 1524:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      exp_reg_1_0 <= exp_reg_0_0; // @[FloatingPointDesigns.scala 1693:22]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1524:28]
      exp_reg_1_1 <= 8'h0; // @[FloatingPointDesigns.scala 1524:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      exp_reg_1_1 <= exp_reg_0_1; // @[FloatingPointDesigns.scala 1693:22]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1524:28]
      exp_reg_2_0 <= 8'h0; // @[FloatingPointDesigns.scala 1524:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      exp_reg_2_0 <= exp_reg_1_0; // @[FloatingPointDesigns.scala 1693:22]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1524:28]
      exp_reg_2_1 <= 8'h0; // @[FloatingPointDesigns.scala 1524:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      exp_reg_2_1 <= exp_reg_1_1; // @[FloatingPointDesigns.scala 1693:22]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1525:28]
      frac_reg_0_0 <= 23'h0; // @[FloatingPointDesigns.scala 1525:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      frac_reg_0_0 <= frac_0; // @[FloatingPointDesigns.scala 1644:19]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1525:28]
      frac_reg_0_1 <= 23'h0; // @[FloatingPointDesigns.scala 1525:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      frac_reg_0_1 <= frac_1; // @[FloatingPointDesigns.scala 1644:19]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1525:28]
      frac_reg_1_0 <= 23'h0; // @[FloatingPointDesigns.scala 1525:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      frac_reg_1_0 <= frac_reg_0_0; // @[FloatingPointDesigns.scala 1694:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1525:28]
      frac_reg_1_1 <= 23'h0; // @[FloatingPointDesigns.scala 1525:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      frac_reg_1_1 <= frac_reg_0_1; // @[FloatingPointDesigns.scala 1694:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1525:28]
      frac_reg_2_0 <= 23'h0; // @[FloatingPointDesigns.scala 1525:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      frac_reg_2_0 <= frac_reg_1_0; // @[FloatingPointDesigns.scala 1694:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1525:28]
      frac_reg_2_1 <= 23'h0; // @[FloatingPointDesigns.scala 1525:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      frac_reg_2_1 <= frac_reg_1_1; // @[FloatingPointDesigns.scala 1694:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1526:28]
      wfrac_reg_0_0 <= 24'h0; // @[FloatingPointDesigns.scala 1526:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      wfrac_reg_0_0 <= whole_frac_0; // @[FloatingPointDesigns.scala 1645:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1526:28]
      wfrac_reg_0_1 <= 24'h0; // @[FloatingPointDesigns.scala 1526:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      wfrac_reg_0_1 <= whole_frac_1; // @[FloatingPointDesigns.scala 1645:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1526:28]
      wfrac_reg_1_0 <= 24'h0; // @[FloatingPointDesigns.scala 1526:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      wfrac_reg_1_0 <= wfrac_reg_0_0; // @[FloatingPointDesigns.scala 1695:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1526:28]
      wfrac_reg_1_1 <= 24'h0; // @[FloatingPointDesigns.scala 1526:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      wfrac_reg_1_1 <= wfrac_reg_0_1; // @[FloatingPointDesigns.scala 1695:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1526:28]
      wfrac_reg_2_0 <= 24'h0; // @[FloatingPointDesigns.scala 1526:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      wfrac_reg_2_0 <= wfrac_reg_1_0; // @[FloatingPointDesigns.scala 1695:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1526:28]
      wfrac_reg_2_1 <= 24'h0; // @[FloatingPointDesigns.scala 1526:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      wfrac_reg_2_1 <= wfrac_reg_1_1; // @[FloatingPointDesigns.scala 1695:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1528:35]
      subber_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1528:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      subber_out_s_reg_0 <= subber_io_out_s; // @[FloatingPointDesigns.scala 1647:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1528:35]
      subber_out_s_reg_1 <= 8'h0; // @[FloatingPointDesigns.scala 1528:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      subber_out_s_reg_1 <= subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1698:31]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1529:35]
      subber_out_c_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1529:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      subber_out_c_reg_0 <= subber_io_out_c; // @[FloatingPointDesigns.scala 1648:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1529:35]
      subber_out_c_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1529:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      subber_out_c_reg_1 <= subber_out_c_reg_0; // @[FloatingPointDesigns.scala 1699:31]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1531:39]
      wire_temp_add_in_reg_0_0 <= 24'h0; // @[FloatingPointDesigns.scala 1531:39]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1581:39]
        wire_temp_add_in_reg_0_0 <= _wire_temp_add_in_0_T; // @[FloatingPointDesigns.scala 1586:27]
      end else begin
        wire_temp_add_in_reg_0_0 <= wfrac_reg_2_0; // @[FloatingPointDesigns.scala 1593:27]
      end
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1531:39]
      wire_temp_add_in_reg_0_1 <= 24'h0; // @[FloatingPointDesigns.scala 1531:39]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1581:39]
        wire_temp_add_in_reg_0_1 <= wfrac_reg_2_1; // @[FloatingPointDesigns.scala 1587:27]
      end else begin
        wire_temp_add_in_reg_0_1 <= _wire_temp_add_in_1_T; // @[FloatingPointDesigns.scala 1594:27]
      end
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1531:39]
      wire_temp_add_in_reg_1_0 <= 24'h0; // @[FloatingPointDesigns.scala 1531:39]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      wire_temp_add_in_reg_1_0 <= wire_temp_add_in_reg_0_0; // @[FloatingPointDesigns.scala 1701:35]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1531:39]
      wire_temp_add_in_reg_1_1 <= 24'h0; // @[FloatingPointDesigns.scala 1531:39]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      wire_temp_add_in_reg_1_1 <= wire_temp_add_in_reg_0_1; // @[FloatingPointDesigns.scala 1701:35]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1533:31]
      ref_s_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1533:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1581:39]
        ref_s_reg_0 <= sign_reg_2_1; // @[FloatingPointDesigns.scala 1584:13]
      end else begin
        ref_s_reg_0 <= sign_reg_2_0; // @[FloatingPointDesigns.scala 1591:13]
      end
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1533:31]
      ref_s_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1533:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_s_reg_1 <= ref_s_reg_0; // @[FloatingPointDesigns.scala 1680:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1533:31]
      ref_s_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1533:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_s_reg_2 <= ref_s_reg_1; // @[FloatingPointDesigns.scala 1680:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1533:31]
      ref_s_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1533:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_s_reg_3 <= ref_s_reg_2; // @[FloatingPointDesigns.scala 1680:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1533:31]
      ref_s_reg_4 <= 1'h0; // @[FloatingPointDesigns.scala 1533:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_s_reg_4 <= ref_s_reg_3; // @[FloatingPointDesigns.scala 1680:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1533:31]
      ref_s_reg_5 <= 1'h0; // @[FloatingPointDesigns.scala 1533:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_s_reg_5 <= ref_s_reg_4; // @[FloatingPointDesigns.scala 1680:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1533:31]
      ref_s_reg_6 <= 1'h0; // @[FloatingPointDesigns.scala 1533:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_s_reg_6 <= ref_s_reg_5; // @[FloatingPointDesigns.scala 1680:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1533:31]
      ref_s_reg_7 <= 1'h0; // @[FloatingPointDesigns.scala 1533:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_s_reg_7 <= ref_s_reg_6; // @[FloatingPointDesigns.scala 1680:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1534:31]
      ref_frac_reg_0 <= 23'h0; // @[FloatingPointDesigns.scala 1534:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1581:39]
        ref_frac_reg_0 <= frac_reg_2_1; // @[FloatingPointDesigns.scala 1585:16]
      end else begin
        ref_frac_reg_0 <= frac_reg_2_0; // @[FloatingPointDesigns.scala 1592:16]
      end
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1534:31]
      ref_frac_reg_1 <= 23'h0; // @[FloatingPointDesigns.scala 1534:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_frac_reg_1 <= ref_frac_reg_0; // @[FloatingPointDesigns.scala 1681:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1534:31]
      ref_frac_reg_2 <= 23'h0; // @[FloatingPointDesigns.scala 1534:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_frac_reg_2 <= ref_frac_reg_1; // @[FloatingPointDesigns.scala 1681:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1534:31]
      ref_frac_reg_3 <= 23'h0; // @[FloatingPointDesigns.scala 1534:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_frac_reg_3 <= ref_frac_reg_2; // @[FloatingPointDesigns.scala 1681:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1534:31]
      ref_frac_reg_4 <= 23'h0; // @[FloatingPointDesigns.scala 1534:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_frac_reg_4 <= ref_frac_reg_3; // @[FloatingPointDesigns.scala 1681:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1534:31]
      ref_frac_reg_5 <= 23'h0; // @[FloatingPointDesigns.scala 1534:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_frac_reg_5 <= ref_frac_reg_4; // @[FloatingPointDesigns.scala 1681:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1534:31]
      ref_frac_reg_6 <= 23'h0; // @[FloatingPointDesigns.scala 1534:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_frac_reg_6 <= ref_frac_reg_5; // @[FloatingPointDesigns.scala 1681:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1534:31]
      ref_frac_reg_7 <= 23'h0; // @[FloatingPointDesigns.scala 1534:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_frac_reg_7 <= ref_frac_reg_6; // @[FloatingPointDesigns.scala 1681:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1535:31]
      ref_exp_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1535:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1581:39]
        ref_exp_reg_0 <= exp_reg_2_1; // @[FloatingPointDesigns.scala 1582:15]
      end else begin
        ref_exp_reg_0 <= exp_reg_2_0; // @[FloatingPointDesigns.scala 1589:15]
      end
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1535:31]
      ref_exp_reg_1 <= 8'h0; // @[FloatingPointDesigns.scala 1535:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_exp_reg_1 <= ref_exp_reg_0; // @[FloatingPointDesigns.scala 1682:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1535:31]
      ref_exp_reg_2 <= 8'h0; // @[FloatingPointDesigns.scala 1535:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_exp_reg_2 <= ref_exp_reg_1; // @[FloatingPointDesigns.scala 1682:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1535:31]
      ref_exp_reg_3 <= 8'h0; // @[FloatingPointDesigns.scala 1535:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_exp_reg_3 <= ref_exp_reg_2; // @[FloatingPointDesigns.scala 1682:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1535:31]
      ref_exp_reg_4 <= 8'h0; // @[FloatingPointDesigns.scala 1535:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_exp_reg_4 <= ref_exp_reg_3; // @[FloatingPointDesigns.scala 1682:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1535:31]
      ref_exp_reg_5 <= 8'h0; // @[FloatingPointDesigns.scala 1535:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_exp_reg_5 <= ref_exp_reg_4; // @[FloatingPointDesigns.scala 1682:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1535:31]
      ref_exp_reg_6 <= 8'h0; // @[FloatingPointDesigns.scala 1535:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_exp_reg_6 <= ref_exp_reg_5; // @[FloatingPointDesigns.scala 1682:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1535:31]
      ref_exp_reg_7 <= 8'h0; // @[FloatingPointDesigns.scala 1535:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      ref_exp_reg_7 <= ref_exp_reg_6; // @[FloatingPointDesigns.scala 1682:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1536:31]
      sub_exp_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1536:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1581:39]
        sub_exp_reg_0 <= cmpl_subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1583:15]
      end else begin
        sub_exp_reg_0 <= subber_out_s_reg_1; // @[FloatingPointDesigns.scala 1590:15]
      end
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1536:31]
      sub_exp_reg_1 <= 8'h0; // @[FloatingPointDesigns.scala 1536:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sub_exp_reg_1 <= sub_exp_reg_0; // @[FloatingPointDesigns.scala 1683:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1536:31]
      sub_exp_reg_2 <= 8'h0; // @[FloatingPointDesigns.scala 1536:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sub_exp_reg_2 <= sub_exp_reg_1; // @[FloatingPointDesigns.scala 1683:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1536:31]
      sub_exp_reg_3 <= 8'h0; // @[FloatingPointDesigns.scala 1536:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sub_exp_reg_3 <= sub_exp_reg_2; // @[FloatingPointDesigns.scala 1683:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1536:31]
      sub_exp_reg_4 <= 8'h0; // @[FloatingPointDesigns.scala 1536:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sub_exp_reg_4 <= sub_exp_reg_3; // @[FloatingPointDesigns.scala 1683:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1536:31]
      sub_exp_reg_5 <= 8'h0; // @[FloatingPointDesigns.scala 1536:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sub_exp_reg_5 <= sub_exp_reg_4; // @[FloatingPointDesigns.scala 1683:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1536:31]
      sub_exp_reg_6 <= 8'h0; // @[FloatingPointDesigns.scala 1536:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sub_exp_reg_6 <= sub_exp_reg_5; // @[FloatingPointDesigns.scala 1683:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1536:31]
      sub_exp_reg_7 <= 8'h0; // @[FloatingPointDesigns.scala 1536:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      sub_exp_reg_7 <= sub_exp_reg_6; // @[FloatingPointDesigns.scala 1683:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1538:37]
      adder_io_out_s_reg_0 <= 24'h0; // @[FloatingPointDesigns.scala 1538:37]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      adder_io_out_s_reg_0 <= adder_io_out_s; // @[FloatingPointDesigns.scala 1663:29]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1538:37]
      adder_io_out_s_reg_1 <= 24'h0; // @[FloatingPointDesigns.scala 1538:37]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      adder_io_out_s_reg_1 <= adder_io_out_s_reg_0; // @[FloatingPointDesigns.scala 1692:33]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1538:37]
      adder_io_out_s_reg_2 <= 24'h0; // @[FloatingPointDesigns.scala 1538:37]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      adder_io_out_s_reg_2 <= adder_io_out_s_reg_1; // @[FloatingPointDesigns.scala 1692:33]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1539:37]
      adder_io_out_c_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1539:37]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      adder_io_out_c_reg_0 <= adder_io_out_c; // @[FloatingPointDesigns.scala 1664:29]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1541:35]
      new_s_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1541:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      new_s_reg_0 <= new_s; // @[FloatingPointDesigns.scala 1657:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1541:35]
      new_s_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1541:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      new_s_reg_1 <= new_s_reg_0; // @[FloatingPointDesigns.scala 1688:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1541:35]
      new_s_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1541:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      new_s_reg_2 <= new_s_reg_1; // @[FloatingPointDesigns.scala 1688:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1541:35]
      new_s_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1541:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      new_s_reg_3 <= new_s_reg_2; // @[FloatingPointDesigns.scala 1688:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1541:35]
      new_s_reg_4 <= 1'h0; // @[FloatingPointDesigns.scala 1541:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      new_s_reg_4 <= new_s_reg_3; // @[FloatingPointDesigns.scala 1688:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1541:35]
      new_s_reg_5 <= 1'h0; // @[FloatingPointDesigns.scala 1541:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1707:20]
      if (io_in_a_reg_10[30:0] == 31'h0 & io_in_b_reg_10[30:0] == 31'h0) begin // @[FloatingPointDesigns.scala 1708:86]
        new_s_reg_5 <= 1'h0; // @[FloatingPointDesigns.scala 1709:22]
      end else if (sub_exp_reg_7 >= 8'h17) begin // @[FloatingPointDesigns.scala 1712:48]
        new_s_reg_5 <= ref_s_reg_7; // @[FloatingPointDesigns.scala 1713:22]
      end else begin
        new_s_reg_5 <= _GEN_154;
      end
    end
    new_out_frac_reg_0 <= _GEN_170[22:0]; // @[FloatingPointDesigns.scala 1542:{35,35}]
    new_out_exp_reg_0 <= _GEN_171[7:0]; // @[FloatingPointDesigns.scala 1543:{35,35}]
    if (reset) begin // @[FloatingPointDesigns.scala 1544:24]
      E_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1544:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      E_reg_0 <= E; // @[FloatingPointDesigns.scala 1660:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1544:24]
      E_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1544:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      E_reg_1 <= E_reg_0; // @[FloatingPointDesigns.scala 1686:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1544:24]
      E_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1544:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      E_reg_2 <= E_reg_1; // @[FloatingPointDesigns.scala 1686:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1544:24]
      E_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1544:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      E_reg_3 <= E_reg_2; // @[FloatingPointDesigns.scala 1686:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1544:24]
      E_reg_4 <= 1'h0; // @[FloatingPointDesigns.scala 1544:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      E_reg_4 <= E_reg_3; // @[FloatingPointDesigns.scala 1686:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1545:24]
      D_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1545:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      D_reg_0 <= D; // @[FloatingPointDesigns.scala 1661:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1545:24]
      D_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1545:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      D_reg_1 <= D_reg_0; // @[FloatingPointDesigns.scala 1687:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1545:24]
      D_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1545:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      D_reg_2 <= D_reg_1; // @[FloatingPointDesigns.scala 1687:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1545:24]
      D_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1545:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      D_reg_3 <= D_reg_2; // @[FloatingPointDesigns.scala 1687:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1545:24]
      D_reg_4 <= 1'h0; // @[FloatingPointDesigns.scala 1545:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      D_reg_4 <= D_reg_3; // @[FloatingPointDesigns.scala 1687:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1547:35]
      adder_result_reg_0 <= 24'h0; // @[FloatingPointDesigns.scala 1547:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      if (new_s_reg_1 & ^_adder_result_T) begin // @[FloatingPointDesigns.scala 1628:24]
        adder_result_reg_0 <= cmpl_adder_io_out_s_reg_0;
      end else begin
        adder_result_reg_0 <= adder_io_out_s_reg_2;
      end
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1547:35]
      adder_result_reg_1 <= 24'h0; // @[FloatingPointDesigns.scala 1547:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      adder_result_reg_1 <= adder_result_reg_0; // @[FloatingPointDesigns.scala 1691:31]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1547:35]
      adder_result_reg_2 <= 24'h0; // @[FloatingPointDesigns.scala 1547:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      adder_result_reg_2 <= adder_result_reg_1; // @[FloatingPointDesigns.scala 1691:31]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1549:33]
      leadingOne_reg_0 <= 6'h0; // @[FloatingPointDesigns.scala 1549:33]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      leadingOne_reg_0 <= leadingOne; // @[FloatingPointDesigns.scala 1668:25]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1549:33]
      leadingOne_reg_1 <= 6'h0; // @[FloatingPointDesigns.scala 1549:33]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      leadingOne_reg_1 <= leadingOne_reg_0; // @[FloatingPointDesigns.scala 1700:29]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1551:30]
      io_in_a_reg_0 <= 32'h0; // @[FloatingPointDesigns.scala 1551:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_a_reg_0 <= io_in_a; // @[FloatingPointDesigns.scala 1639:22]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1551:30]
      io_in_a_reg_1 <= 32'h0; // @[FloatingPointDesigns.scala 1551:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_a_reg_1 <= io_in_a_reg_0; // @[FloatingPointDesigns.scala 1676:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1551:30]
      io_in_a_reg_2 <= 32'h0; // @[FloatingPointDesigns.scala 1551:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_a_reg_2 <= io_in_a_reg_1; // @[FloatingPointDesigns.scala 1676:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1551:30]
      io_in_a_reg_3 <= 32'h0; // @[FloatingPointDesigns.scala 1551:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_a_reg_3 <= io_in_a_reg_2; // @[FloatingPointDesigns.scala 1676:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1551:30]
      io_in_a_reg_4 <= 32'h0; // @[FloatingPointDesigns.scala 1551:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_a_reg_4 <= io_in_a_reg_3; // @[FloatingPointDesigns.scala 1676:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1551:30]
      io_in_a_reg_5 <= 32'h0; // @[FloatingPointDesigns.scala 1551:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_a_reg_5 <= io_in_a_reg_4; // @[FloatingPointDesigns.scala 1676:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1551:30]
      io_in_a_reg_6 <= 32'h0; // @[FloatingPointDesigns.scala 1551:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_a_reg_6 <= io_in_a_reg_5; // @[FloatingPointDesigns.scala 1676:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1551:30]
      io_in_a_reg_7 <= 32'h0; // @[FloatingPointDesigns.scala 1551:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_a_reg_7 <= io_in_a_reg_6; // @[FloatingPointDesigns.scala 1676:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1551:30]
      io_in_a_reg_8 <= 32'h0; // @[FloatingPointDesigns.scala 1551:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_a_reg_8 <= io_in_a_reg_7; // @[FloatingPointDesigns.scala 1676:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1551:30]
      io_in_a_reg_9 <= 32'h0; // @[FloatingPointDesigns.scala 1551:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_a_reg_9 <= io_in_a_reg_8; // @[FloatingPointDesigns.scala 1676:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1551:30]
      io_in_a_reg_10 <= 32'h0; // @[FloatingPointDesigns.scala 1551:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_a_reg_10 <= io_in_a_reg_9; // @[FloatingPointDesigns.scala 1676:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1552:30]
      io_in_b_reg_0 <= 32'h0; // @[FloatingPointDesigns.scala 1552:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_b_reg_0 <= io_in_b; // @[FloatingPointDesigns.scala 1640:22]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1552:30]
      io_in_b_reg_1 <= 32'h0; // @[FloatingPointDesigns.scala 1552:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_b_reg_1 <= io_in_b_reg_0; // @[FloatingPointDesigns.scala 1677:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1552:30]
      io_in_b_reg_2 <= 32'h0; // @[FloatingPointDesigns.scala 1552:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_b_reg_2 <= io_in_b_reg_1; // @[FloatingPointDesigns.scala 1677:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1552:30]
      io_in_b_reg_3 <= 32'h0; // @[FloatingPointDesigns.scala 1552:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_b_reg_3 <= io_in_b_reg_2; // @[FloatingPointDesigns.scala 1677:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1552:30]
      io_in_b_reg_4 <= 32'h0; // @[FloatingPointDesigns.scala 1552:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_b_reg_4 <= io_in_b_reg_3; // @[FloatingPointDesigns.scala 1677:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1552:30]
      io_in_b_reg_5 <= 32'h0; // @[FloatingPointDesigns.scala 1552:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_b_reg_5 <= io_in_b_reg_4; // @[FloatingPointDesigns.scala 1677:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1552:30]
      io_in_b_reg_6 <= 32'h0; // @[FloatingPointDesigns.scala 1552:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_b_reg_6 <= io_in_b_reg_5; // @[FloatingPointDesigns.scala 1677:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1552:30]
      io_in_b_reg_7 <= 32'h0; // @[FloatingPointDesigns.scala 1552:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_b_reg_7 <= io_in_b_reg_6; // @[FloatingPointDesigns.scala 1677:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1552:30]
      io_in_b_reg_8 <= 32'h0; // @[FloatingPointDesigns.scala 1552:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_b_reg_8 <= io_in_b_reg_7; // @[FloatingPointDesigns.scala 1677:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1552:30]
      io_in_b_reg_9 <= 32'h0; // @[FloatingPointDesigns.scala 1552:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_b_reg_9 <= io_in_b_reg_8; // @[FloatingPointDesigns.scala 1677:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1552:30]
      io_in_b_reg_10 <= 32'h0; // @[FloatingPointDesigns.scala 1552:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      io_in_b_reg_10 <= io_in_b_reg_9; // @[FloatingPointDesigns.scala 1677:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1554:36]
      subber2_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1554:36]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      subber2_out_s_reg_0 <= subber2_io_out_s; // @[FloatingPointDesigns.scala 1670:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1555:36]
      subber2_out_c_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1555:36]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1638:19]
      subber2_out_c_reg_0 <= subber2_io_out_c; // @[FloatingPointDesigns.scala 1671:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1576:40]
      cmpl_subber_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1576:40]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1577:19]
      cmpl_subber_out_s_reg_0 <= _cmpl_subber_out_s_reg_0_T_2; // @[FloatingPointDesigns.scala 1578:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1597:44]
      cmpl_wire_temp_add_in_reg_0_0 <= 24'h0; // @[FloatingPointDesigns.scala 1597:44]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1598:19]
      cmpl_wire_temp_add_in_reg_0_0 <= _cmpl_wire_temp_add_in_reg_0_0_T_2; // @[FloatingPointDesigns.scala 1599:39]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1597:44]
      cmpl_wire_temp_add_in_reg_0_1 <= 24'h0; // @[FloatingPointDesigns.scala 1597:44]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1598:19]
      cmpl_wire_temp_add_in_reg_0_1 <= _cmpl_wire_temp_add_in_reg_0_1_T_2; // @[FloatingPointDesigns.scala 1600:39]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1621:42]
      cmpl_adder_io_out_s_reg_0 <= 24'h0; // @[FloatingPointDesigns.scala 1621:42]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1623:19]
      cmpl_adder_io_out_s_reg_0 <= _cmpl_adder_io_out_s_reg_0_T_2; // @[FloatingPointDesigns.scala 1624:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1705:28]
      reg_out_s <= 32'h0; // @[FloatingPointDesigns.scala 1705:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1707:20]
      reg_out_s <= _reg_out_s_T_1; // @[FloatingPointDesigns.scala 1744:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sign_reg_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sign_reg_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sign_reg_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  sign_reg_1_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  sign_reg_2_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  sign_reg_2_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  sign_reg_3_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  sign_reg_3_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sign_reg_4_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sign_reg_4_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  sign_reg_5_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  sign_reg_5_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  sign_reg_6_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  sign_reg_6_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  sign_reg_7_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  sign_reg_7_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  sign_reg_8_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  sign_reg_8_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  sign_reg_9_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sign_reg_9_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  sign_reg_10_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  sign_reg_10_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  exp_reg_0_0 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  exp_reg_0_1 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  exp_reg_1_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  exp_reg_1_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  exp_reg_2_0 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  exp_reg_2_1 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  frac_reg_0_0 = _RAND_28[22:0];
  _RAND_29 = {1{`RANDOM}};
  frac_reg_0_1 = _RAND_29[22:0];
  _RAND_30 = {1{`RANDOM}};
  frac_reg_1_0 = _RAND_30[22:0];
  _RAND_31 = {1{`RANDOM}};
  frac_reg_1_1 = _RAND_31[22:0];
  _RAND_32 = {1{`RANDOM}};
  frac_reg_2_0 = _RAND_32[22:0];
  _RAND_33 = {1{`RANDOM}};
  frac_reg_2_1 = _RAND_33[22:0];
  _RAND_34 = {1{`RANDOM}};
  wfrac_reg_0_0 = _RAND_34[23:0];
  _RAND_35 = {1{`RANDOM}};
  wfrac_reg_0_1 = _RAND_35[23:0];
  _RAND_36 = {1{`RANDOM}};
  wfrac_reg_1_0 = _RAND_36[23:0];
  _RAND_37 = {1{`RANDOM}};
  wfrac_reg_1_1 = _RAND_37[23:0];
  _RAND_38 = {1{`RANDOM}};
  wfrac_reg_2_0 = _RAND_38[23:0];
  _RAND_39 = {1{`RANDOM}};
  wfrac_reg_2_1 = _RAND_39[23:0];
  _RAND_40 = {1{`RANDOM}};
  subber_out_s_reg_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  subber_out_s_reg_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  subber_out_c_reg_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  subber_out_c_reg_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  wire_temp_add_in_reg_0_0 = _RAND_44[23:0];
  _RAND_45 = {1{`RANDOM}};
  wire_temp_add_in_reg_0_1 = _RAND_45[23:0];
  _RAND_46 = {1{`RANDOM}};
  wire_temp_add_in_reg_1_0 = _RAND_46[23:0];
  _RAND_47 = {1{`RANDOM}};
  wire_temp_add_in_reg_1_1 = _RAND_47[23:0];
  _RAND_48 = {1{`RANDOM}};
  ref_s_reg_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  ref_s_reg_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  ref_s_reg_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  ref_s_reg_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  ref_s_reg_4 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  ref_s_reg_5 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  ref_s_reg_6 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  ref_s_reg_7 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  ref_frac_reg_0 = _RAND_56[22:0];
  _RAND_57 = {1{`RANDOM}};
  ref_frac_reg_1 = _RAND_57[22:0];
  _RAND_58 = {1{`RANDOM}};
  ref_frac_reg_2 = _RAND_58[22:0];
  _RAND_59 = {1{`RANDOM}};
  ref_frac_reg_3 = _RAND_59[22:0];
  _RAND_60 = {1{`RANDOM}};
  ref_frac_reg_4 = _RAND_60[22:0];
  _RAND_61 = {1{`RANDOM}};
  ref_frac_reg_5 = _RAND_61[22:0];
  _RAND_62 = {1{`RANDOM}};
  ref_frac_reg_6 = _RAND_62[22:0];
  _RAND_63 = {1{`RANDOM}};
  ref_frac_reg_7 = _RAND_63[22:0];
  _RAND_64 = {1{`RANDOM}};
  ref_exp_reg_0 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  ref_exp_reg_1 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  ref_exp_reg_2 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  ref_exp_reg_3 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  ref_exp_reg_4 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  ref_exp_reg_5 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  ref_exp_reg_6 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  ref_exp_reg_7 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  sub_exp_reg_0 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  sub_exp_reg_1 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  sub_exp_reg_2 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  sub_exp_reg_3 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  sub_exp_reg_4 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  sub_exp_reg_5 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  sub_exp_reg_6 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  sub_exp_reg_7 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  adder_io_out_s_reg_0 = _RAND_80[23:0];
  _RAND_81 = {1{`RANDOM}};
  adder_io_out_s_reg_1 = _RAND_81[23:0];
  _RAND_82 = {1{`RANDOM}};
  adder_io_out_s_reg_2 = _RAND_82[23:0];
  _RAND_83 = {1{`RANDOM}};
  adder_io_out_c_reg_0 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  new_s_reg_0 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  new_s_reg_1 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  new_s_reg_2 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  new_s_reg_3 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  new_s_reg_4 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  new_s_reg_5 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  new_out_frac_reg_0 = _RAND_90[22:0];
  _RAND_91 = {1{`RANDOM}};
  new_out_exp_reg_0 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  E_reg_0 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  E_reg_1 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  E_reg_2 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  E_reg_3 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  E_reg_4 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  D_reg_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  D_reg_1 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  D_reg_2 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  D_reg_3 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  D_reg_4 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  adder_result_reg_0 = _RAND_102[23:0];
  _RAND_103 = {1{`RANDOM}};
  adder_result_reg_1 = _RAND_103[23:0];
  _RAND_104 = {1{`RANDOM}};
  adder_result_reg_2 = _RAND_104[23:0];
  _RAND_105 = {1{`RANDOM}};
  leadingOne_reg_0 = _RAND_105[5:0];
  _RAND_106 = {1{`RANDOM}};
  leadingOne_reg_1 = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  io_in_a_reg_0 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  io_in_a_reg_1 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  io_in_a_reg_2 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  io_in_a_reg_3 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  io_in_a_reg_4 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  io_in_a_reg_5 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  io_in_a_reg_6 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  io_in_a_reg_7 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  io_in_a_reg_8 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  io_in_a_reg_9 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  io_in_a_reg_10 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  io_in_b_reg_0 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  io_in_b_reg_1 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  io_in_b_reg_2 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  io_in_b_reg_3 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  io_in_b_reg_4 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  io_in_b_reg_5 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  io_in_b_reg_6 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  io_in_b_reg_7 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  io_in_b_reg_8 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  io_in_b_reg_9 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  io_in_b_reg_10 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  subber2_out_s_reg_0 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  subber2_out_c_reg_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  cmpl_subber_out_s_reg_0 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  cmpl_wire_temp_add_in_reg_0_0 = _RAND_132[23:0];
  _RAND_133 = {1{`RANDOM}};
  cmpl_wire_temp_add_in_reg_0_1 = _RAND_133[23:0];
  _RAND_134 = {1{`RANDOM}};
  cmpl_adder_io_out_s_reg_0 = _RAND_134[23:0];
  _RAND_135 = {1{`RANDOM}};
  reg_out_s = _RAND_135[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FP_subtractor_13ccs(
  input         clock,
  input         reset,
  input         io_in_en,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
  wire  FP_adder_clock; // @[FloatingPointDesigns.scala 1759:26]
  wire  FP_adder_reset; // @[FloatingPointDesigns.scala 1759:26]
  wire  FP_adder_io_in_en; // @[FloatingPointDesigns.scala 1759:26]
  wire [31:0] FP_adder_io_in_a; // @[FloatingPointDesigns.scala 1759:26]
  wire [31:0] FP_adder_io_in_b; // @[FloatingPointDesigns.scala 1759:26]
  wire [31:0] FP_adder_io_out_s; // @[FloatingPointDesigns.scala 1759:26]
  wire  _adjusted_in_b_T_1 = ~io_in_b[31]; // @[FloatingPointDesigns.scala 1762:23]
  FP_adder_13ccs FP_adder ( // @[FloatingPointDesigns.scala 1759:26]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_en(FP_adder_io_in_en),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  assign io_out_s = FP_adder_io_out_s; // @[FloatingPointDesigns.scala 1766:14]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1763:23]
  assign FP_adder_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 1764:22]
  assign FP_adder_io_in_b = {_adjusted_in_b_T_1,io_in_b[30:0]}; // @[FloatingPointDesigns.scala 1762:41]
endmodule
module multiplier(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [47:0] io_out_s
);
  assign io_out_s = io_in_a * io_in_b; // @[BinaryDesigns.scala 81:23]
endmodule
module twoscomplement(
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _x_T = ~io_in; // @[BinaryDesigns.scala 25:16]
  assign io_out = 8'h1 + _x_T; // @[BinaryDesigns.scala 25:14]
endmodule
module full_adder_2(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s,
  output       io_out_c
);
  wire [8:0] _result_T = io_in_a + io_in_b; // @[BinaryDesigns.scala 55:23]
  wire [9:0] _result_T_1 = {{1'd0}, _result_T}; // @[BinaryDesigns.scala 55:34]
  wire [8:0] result = _result_T_1[8:0]; // @[BinaryDesigns.scala 54:22 55:12]
  assign io_out_s = result[7:0]; // @[BinaryDesigns.scala 56:23]
  assign io_out_c = result[8]; // @[BinaryDesigns.scala 57:23]
endmodule
module FP_multiplier_10ccs(
  input         clock,
  input         reset,
  input         io_in_en,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
`endif // RANDOMIZE_REG_INIT
  wire [23:0] multiplier_io_in_a; // @[FloatingPointDesigns.scala 1830:28]
  wire [23:0] multiplier_io_in_b; // @[FloatingPointDesigns.scala 1830:28]
  wire [47:0] multiplier_io_out_s; // @[FloatingPointDesigns.scala 1830:28]
  wire [7:0] subber_io_in_a; // @[FloatingPointDesigns.scala 1837:24]
  wire [7:0] subber_io_in_b; // @[FloatingPointDesigns.scala 1837:24]
  wire [7:0] subber_io_out_s; // @[FloatingPointDesigns.scala 1837:24]
  wire  subber_io_out_c; // @[FloatingPointDesigns.scala 1837:24]
  wire [7:0] complementN_io_in; // @[FloatingPointDesigns.scala 1846:29]
  wire [7:0] complementN_io_out; // @[FloatingPointDesigns.scala 1846:29]
  wire [7:0] adderN_io_in_a; // @[FloatingPointDesigns.scala 1863:24]
  wire [7:0] adderN_io_in_b; // @[FloatingPointDesigns.scala 1863:24]
  wire [7:0] adderN_io_out_s; // @[FloatingPointDesigns.scala 1863:24]
  wire  adderN_io_out_c; // @[FloatingPointDesigns.scala 1863:24]
  wire  s_0 = io_in_a[31]; // @[FloatingPointDesigns.scala 1796:20]
  wire  s_1 = io_in_b[31]; // @[FloatingPointDesigns.scala 1797:20]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FloatingPointDesigns.scala 1801:64]
  wire [8:0] _GEN_63 = {{1'd0}, io_in_a[30:23]}; // @[FloatingPointDesigns.scala 1801:36]
  wire [7:0] _GEN_0 = io_in_a[30:23] < 8'h1 ? 8'h1 : io_in_a[30:23]; // @[FloatingPointDesigns.scala 1803:45 1804:14 1806:14]
  wire [8:0] _GEN_1 = _GEN_63 > _T_2 ? _T_2 : {{1'd0}, _GEN_0}; // @[FloatingPointDesigns.scala 1801:71 1802:14]
  wire [8:0] _GEN_64 = {{1'd0}, io_in_b[30:23]}; // @[FloatingPointDesigns.scala 1808:36]
  wire [7:0] _GEN_2 = io_in_b[30:23] < 8'h1 ? 8'h1 : io_in_b[30:23]; // @[FloatingPointDesigns.scala 1810:45 1811:14 1813:14]
  wire [8:0] _GEN_3 = _GEN_64 > _T_2 ? _T_2 : {{1'd0}, _GEN_2}; // @[FloatingPointDesigns.scala 1808:71 1809:14]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FloatingPointDesigns.scala 1818:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FloatingPointDesigns.scala 1819:23]
  wire [23:0] new_frac_0 = {1'h1,frac_0}; // @[FloatingPointDesigns.scala 1823:24]
  wire [23:0] new_frac_1 = {1'h1,frac_1}; // @[FloatingPointDesigns.scala 1824:24]
  reg  s_reg_0_0; // @[FloatingPointDesigns.scala 1826:24]
  reg  s_reg_0_1; // @[FloatingPointDesigns.scala 1826:24]
  reg  s_reg_1_0; // @[FloatingPointDesigns.scala 1826:24]
  reg  s_reg_1_1; // @[FloatingPointDesigns.scala 1826:24]
  reg  s_reg_2_0; // @[FloatingPointDesigns.scala 1826:24]
  reg  s_reg_2_1; // @[FloatingPointDesigns.scala 1826:24]
  reg  s_reg_3_0; // @[FloatingPointDesigns.scala 1826:24]
  reg  s_reg_3_1; // @[FloatingPointDesigns.scala 1826:24]
  reg  s_reg_4_0; // @[FloatingPointDesigns.scala 1826:24]
  reg  s_reg_4_1; // @[FloatingPointDesigns.scala 1826:24]
  reg [7:0] exp_reg_0_0; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_0_1; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_1_0; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_1_1; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_2_0; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_2_1; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_3_0; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_3_1; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_4_0; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_4_1; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_5_0; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_5_1; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_6_0; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_6_1; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_7_0; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_7_1; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_8_0; // @[FloatingPointDesigns.scala 1827:26]
  reg [7:0] exp_reg_8_1; // @[FloatingPointDesigns.scala 1827:26]
  reg [23:0] new_frac_reg_0_0; // @[FloatingPointDesigns.scala 1828:31]
  reg [23:0] new_frac_reg_0_1; // @[FloatingPointDesigns.scala 1828:31]
  reg [23:0] new_frac_reg_1_0; // @[FloatingPointDesigns.scala 1828:31]
  reg [23:0] new_frac_reg_1_1; // @[FloatingPointDesigns.scala 1828:31]
  reg [47:0] multipplier_out_s_reg_0; // @[FloatingPointDesigns.scala 1834:40]
  reg [47:0] multipplier_out_s_reg_1; // @[FloatingPointDesigns.scala 1834:40]
  reg [47:0] multipplier_out_s_reg_2; // @[FloatingPointDesigns.scala 1834:40]
  reg [47:0] multipplier_out_s_reg_3; // @[FloatingPointDesigns.scala 1834:40]
  reg [47:0] multipplier_out_s_reg_4; // @[FloatingPointDesigns.scala 1834:40]
  reg [47:0] multipplier_out_s_reg_5; // @[FloatingPointDesigns.scala 1834:40]
  reg [7:0] subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1842:35]
  reg [7:0] complementN_out_reg_0; // @[FloatingPointDesigns.scala 1849:38]
  reg [7:0] complementN_out_reg_1; // @[FloatingPointDesigns.scala 1849:38]
  reg [7:0] complementN_out_reg_2; // @[FloatingPointDesigns.scala 1849:38]
  wire  new_s = s_reg_4_0 ^ s_reg_4_1; // @[FloatingPointDesigns.scala 1852:26]
  reg  new_s_reg_0; // @[FloatingPointDesigns.scala 1854:28]
  reg  new_s_reg_1; // @[FloatingPointDesigns.scala 1854:28]
  reg  new_s_reg_2; // @[FloatingPointDesigns.scala 1854:28]
  reg  new_s_reg_3; // @[FloatingPointDesigns.scala 1854:28]
  wire  is_exp1_neg_wire = exp_reg_5_1 < 8'h7f; // @[FloatingPointDesigns.scala 1857:40]
  reg  is_exp1_neg_reg_0; // @[FloatingPointDesigns.scala 1859:34]
  reg  is_exp1_neg_reg_1; // @[FloatingPointDesigns.scala 1859:34]
  wire [7:0] _adderN_io_in_a_T_1 = exp_reg_6_0 + 8'h1; // @[FloatingPointDesigns.scala 1867:39]
  reg [7:0] adderN_out_s_reg_0; // @[FloatingPointDesigns.scala 1874:35]
  reg  adderN_out_c_reg_0; // @[FloatingPointDesigns.scala 1875:35]
  reg [7:0] new_exp_reg_0; // @[FloatingPointDesigns.scala 1877:30]
  reg [22:0] new_mant_reg_0; // @[FloatingPointDesigns.scala 1878:31]
  reg [31:0] reg_out_s; // @[FloatingPointDesigns.scala 1880:28]
  wire  _new_exp_reg_0_T_1 = ~adderN_out_c_reg_0; // @[FloatingPointDesigns.scala 1884:55]
  wire [7:0] _new_exp_reg_0_T_2 = ~adderN_out_c_reg_0 ? 8'h1 : adderN_out_s_reg_0; // @[FloatingPointDesigns.scala 1884:54]
  wire  _new_exp_reg_0_T_5 = adderN_out_c_reg_0 | adderN_out_s_reg_0 > 8'hfe; // @[FloatingPointDesigns.scala 1884:142]
  wire [7:0] _new_exp_reg_0_T_6 = adderN_out_c_reg_0 | adderN_out_s_reg_0 > 8'hfe ? 8'hfe : adderN_out_s_reg_0; // @[FloatingPointDesigns.scala 1884:114]
  wire [7:0] _new_exp_reg_0_T_7 = is_exp1_neg_reg_1 ? _new_exp_reg_0_T_2 : _new_exp_reg_0_T_6; // @[FloatingPointDesigns.scala 1884:30]
  wire [22:0] _new_mant_reg_0_T_3 = _new_exp_reg_0_T_1 ? 23'h0 : multipplier_out_s_reg_5[46:24]; // @[FloatingPointDesigns.scala 1885:55]
  wire [22:0] _new_mant_reg_0_T_8 = _new_exp_reg_0_T_5 ? 23'h7fffff : multipplier_out_s_reg_5[46:24]; // @[FloatingPointDesigns.scala 1885:160]
  wire [22:0] _new_mant_reg_0_T_13 = _new_exp_reg_0_T_1 ? 23'h0 : multipplier_out_s_reg_5[45:23]; // @[FloatingPointDesigns.scala 1888:55]
  wire [22:0] _new_mant_reg_0_T_18 = _new_exp_reg_0_T_5 ? 23'h7fffff : multipplier_out_s_reg_5[45:23]; // @[FloatingPointDesigns.scala 1888:156]
  wire [31:0] _reg_out_s_T_1 = {new_s_reg_3,new_exp_reg_0,new_mant_reg_0}; // @[FloatingPointDesigns.scala 1926:53]
  wire [7:0] exp_0 = _GEN_1[7:0]; // @[FloatingPointDesigns.scala 1800:19]
  wire [7:0] exp_1 = _GEN_3[7:0]; // @[FloatingPointDesigns.scala 1800:19]
  multiplier multiplier ( // @[FloatingPointDesigns.scala 1830:28]
    .io_in_a(multiplier_io_in_a),
    .io_in_b(multiplier_io_in_b),
    .io_out_s(multiplier_io_out_s)
  );
  full_subber subber ( // @[FloatingPointDesigns.scala 1837:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  twoscomplement complementN ( // @[FloatingPointDesigns.scala 1846:29]
    .io_in(complementN_io_in),
    .io_out(complementN_io_out)
  );
  full_adder_2 adderN ( // @[FloatingPointDesigns.scala 1863:24]
    .io_in_a(adderN_io_in_a),
    .io_in_b(adderN_io_in_b),
    .io_out_s(adderN_io_out_s),
    .io_out_c(adderN_io_out_c)
  );
  assign io_out_s = reg_out_s; // @[FloatingPointDesigns.scala 1929:14]
  assign multiplier_io_in_a = new_frac_reg_1_0; // @[FloatingPointDesigns.scala 1831:24]
  assign multiplier_io_in_b = new_frac_reg_1_1; // @[FloatingPointDesigns.scala 1832:24]
  assign subber_io_in_a = 8'h7f; // @[FloatingPointDesigns.scala 1838:20]
  assign subber_io_in_b = exp_reg_2_1; // @[FloatingPointDesigns.scala 1839:20]
  assign complementN_io_in = subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1847:23]
  assign adderN_io_in_a = multipplier_out_s_reg_4[47] ? _adderN_io_in_a_T_1 : exp_reg_6_0; // @[FloatingPointDesigns.scala 1866:70 1867:22 1870:22]
  assign adderN_io_in_b = complementN_out_reg_2; // @[FloatingPointDesigns.scala 1866:70 1868:22 1871:22]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 1826:24]
      s_reg_0_0 <= 1'h0; // @[FloatingPointDesigns.scala 1826:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      s_reg_0_0 <= s_0; // @[FloatingPointDesigns.scala 1891:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1826:24]
      s_reg_0_1 <= 1'h0; // @[FloatingPointDesigns.scala 1826:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      s_reg_0_1 <= s_1; // @[FloatingPointDesigns.scala 1891:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1826:24]
      s_reg_1_0 <= 1'h0; // @[FloatingPointDesigns.scala 1826:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      s_reg_1_0 <= s_reg_0_0; // @[FloatingPointDesigns.scala 1908:22]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1826:24]
      s_reg_1_1 <= 1'h0; // @[FloatingPointDesigns.scala 1826:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      s_reg_1_1 <= s_reg_0_1; // @[FloatingPointDesigns.scala 1908:22]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1826:24]
      s_reg_2_0 <= 1'h0; // @[FloatingPointDesigns.scala 1826:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      s_reg_2_0 <= s_reg_1_0; // @[FloatingPointDesigns.scala 1908:22]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1826:24]
      s_reg_2_1 <= 1'h0; // @[FloatingPointDesigns.scala 1826:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      s_reg_2_1 <= s_reg_1_1; // @[FloatingPointDesigns.scala 1908:22]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1826:24]
      s_reg_3_0 <= 1'h0; // @[FloatingPointDesigns.scala 1826:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      s_reg_3_0 <= s_reg_2_0; // @[FloatingPointDesigns.scala 1908:22]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1826:24]
      s_reg_3_1 <= 1'h0; // @[FloatingPointDesigns.scala 1826:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      s_reg_3_1 <= s_reg_2_1; // @[FloatingPointDesigns.scala 1908:22]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1826:24]
      s_reg_4_0 <= 1'h0; // @[FloatingPointDesigns.scala 1826:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      s_reg_4_0 <= s_reg_3_0; // @[FloatingPointDesigns.scala 1908:22]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1826:24]
      s_reg_4_1 <= 1'h0; // @[FloatingPointDesigns.scala 1826:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      s_reg_4_1 <= s_reg_3_1; // @[FloatingPointDesigns.scala 1908:22]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_0_0 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_0_0 <= exp_0; // @[FloatingPointDesigns.scala 1892:18]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_0_1 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_0_1 <= exp_1; // @[FloatingPointDesigns.scala 1892:18]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_1_0 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_1_0 <= exp_reg_0_0; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_1_1 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_1_1 <= exp_reg_0_1; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_2_0 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_2_0 <= exp_reg_1_0; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_2_1 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_2_1 <= exp_reg_1_1; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_3_0 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_3_0 <= exp_reg_2_0; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_3_1 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_3_1 <= exp_reg_2_1; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_4_0 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_4_0 <= exp_reg_3_0; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_4_1 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_4_1 <= exp_reg_3_1; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_5_0 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_5_0 <= exp_reg_4_0; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_5_1 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_5_1 <= exp_reg_4_1; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_6_0 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_6_0 <= exp_reg_5_0; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_6_1 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_6_1 <= exp_reg_5_1; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_7_0 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_7_0 <= exp_reg_6_0; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_7_1 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_7_1 <= exp_reg_6_1; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_8_0 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_8_0 <= exp_reg_7_0; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1827:26]
      exp_reg_8_1 <= 8'h0; // @[FloatingPointDesigns.scala 1827:26]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      exp_reg_8_1 <= exp_reg_7_1; // @[FloatingPointDesigns.scala 1904:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1828:31]
      new_frac_reg_0_0 <= 24'h0; // @[FloatingPointDesigns.scala 1828:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      new_frac_reg_0_0 <= new_frac_0; // @[FloatingPointDesigns.scala 1893:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1828:31]
      new_frac_reg_0_1 <= 24'h0; // @[FloatingPointDesigns.scala 1828:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      new_frac_reg_0_1 <= new_frac_1; // @[FloatingPointDesigns.scala 1893:23]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1828:31]
      new_frac_reg_1_0 <= 24'h0; // @[FloatingPointDesigns.scala 1828:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      new_frac_reg_1_0 <= new_frac_reg_0_0; // @[FloatingPointDesigns.scala 1914:35]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1828:31]
      new_frac_reg_1_1 <= 24'h0; // @[FloatingPointDesigns.scala 1828:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      new_frac_reg_1_1 <= new_frac_reg_0_1; // @[FloatingPointDesigns.scala 1914:35]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1834:40]
      multipplier_out_s_reg_0 <= 48'h0; // @[FloatingPointDesigns.scala 1834:40]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      multipplier_out_s_reg_0 <= multiplier_io_out_s; // @[FloatingPointDesigns.scala 1894:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1834:40]
      multipplier_out_s_reg_1 <= 48'h0; // @[FloatingPointDesigns.scala 1834:40]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      multipplier_out_s_reg_1 <= multipplier_out_s_reg_0; // @[FloatingPointDesigns.scala 1906:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1834:40]
      multipplier_out_s_reg_2 <= 48'h0; // @[FloatingPointDesigns.scala 1834:40]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      multipplier_out_s_reg_2 <= multipplier_out_s_reg_1; // @[FloatingPointDesigns.scala 1906:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1834:40]
      multipplier_out_s_reg_3 <= 48'h0; // @[FloatingPointDesigns.scala 1834:40]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      multipplier_out_s_reg_3 <= multipplier_out_s_reg_2; // @[FloatingPointDesigns.scala 1906:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1834:40]
      multipplier_out_s_reg_4 <= 48'h0; // @[FloatingPointDesigns.scala 1834:40]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      multipplier_out_s_reg_4 <= multipplier_out_s_reg_3; // @[FloatingPointDesigns.scala 1906:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1834:40]
      multipplier_out_s_reg_5 <= 48'h0; // @[FloatingPointDesigns.scala 1834:40]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      multipplier_out_s_reg_5 <= multipplier_out_s_reg_4; // @[FloatingPointDesigns.scala 1906:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1842:35]
      subber_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1842:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      subber_out_s_reg_0 <= subber_io_out_s; // @[FloatingPointDesigns.scala 1895:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1849:38]
      complementN_out_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1849:38]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      complementN_out_reg_0 <= complementN_io_out; // @[FloatingPointDesigns.scala 1897:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1849:38]
      complementN_out_reg_1 <= 8'h0; // @[FloatingPointDesigns.scala 1849:38]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      complementN_out_reg_1 <= complementN_out_reg_0; // @[FloatingPointDesigns.scala 1912:40]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1849:38]
      complementN_out_reg_2 <= 8'h0; // @[FloatingPointDesigns.scala 1849:38]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      complementN_out_reg_2 <= complementN_out_reg_1; // @[FloatingPointDesigns.scala 1912:40]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1854:28]
      new_s_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1854:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      new_s_reg_0 <= new_s; // @[FloatingPointDesigns.scala 1898:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1854:28]
      new_s_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1854:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      new_s_reg_1 <= new_s_reg_0; // @[FloatingPointDesigns.scala 1910:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1854:28]
      new_s_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1854:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      new_s_reg_2 <= new_s_reg_1; // @[FloatingPointDesigns.scala 1910:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1854:28]
      new_s_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1854:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      new_s_reg_3 <= new_s_reg_2; // @[FloatingPointDesigns.scala 1910:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1859:34]
      is_exp1_neg_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1859:34]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      is_exp1_neg_reg_0 <= is_exp1_neg_wire; // @[FloatingPointDesigns.scala 1899:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1859:34]
      is_exp1_neg_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1859:34]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      is_exp1_neg_reg_1 <= is_exp1_neg_reg_0; // @[FloatingPointDesigns.scala 1915:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:35]
      adderN_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1874:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      adderN_out_s_reg_0 <= adderN_io_out_s; // @[FloatingPointDesigns.scala 1900:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:35]
      adderN_out_c_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1875:35]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      adderN_out_c_reg_0 <= adderN_io_out_c; // @[FloatingPointDesigns.scala 1901:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1877:30]
      new_exp_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1877:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      if (multipplier_out_s_reg_5[47]) begin // @[FloatingPointDesigns.scala 1883:72]
        new_exp_reg_0 <= _new_exp_reg_0_T_7; // @[FloatingPointDesigns.scala 1884:24]
      end else begin
        new_exp_reg_0 <= _new_exp_reg_0_T_7; // @[FloatingPointDesigns.scala 1887:24]
      end
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1878:31]
      new_mant_reg_0 <= 23'h0; // @[FloatingPointDesigns.scala 1878:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      if (multipplier_out_s_reg_5[47]) begin // @[FloatingPointDesigns.scala 1883:72]
        if (is_exp1_neg_reg_1) begin // @[FloatingPointDesigns.scala 1885:31]
          new_mant_reg_0 <= _new_mant_reg_0_T_3;
        end else begin
          new_mant_reg_0 <= _new_mant_reg_0_T_8;
        end
      end else if (is_exp1_neg_reg_1) begin // @[FloatingPointDesigns.scala 1888:31]
        new_mant_reg_0 <= _new_mant_reg_0_T_13;
      end else begin
        new_mant_reg_0 <= _new_mant_reg_0_T_18;
      end
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1880:28]
      reg_out_s <= 32'h0; // @[FloatingPointDesigns.scala 1880:28]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1882:19]
      if (exp_reg_8_0 == 8'h0 | exp_reg_8_1 == 8'h0) begin // @[FloatingPointDesigns.scala 1923:60]
        reg_out_s <= 32'h0; // @[FloatingPointDesigns.scala 1924:19]
      end else begin
        reg_out_s <= _reg_out_s_T_1; // @[FloatingPointDesigns.scala 1926:19]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s_reg_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s_reg_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s_reg_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  s_reg_1_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  s_reg_2_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  s_reg_2_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  s_reg_3_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s_reg_3_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  s_reg_4_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  s_reg_4_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  exp_reg_0_0 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  exp_reg_0_1 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  exp_reg_1_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  exp_reg_1_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  exp_reg_2_0 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  exp_reg_2_1 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  exp_reg_3_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  exp_reg_3_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  exp_reg_4_0 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  exp_reg_4_1 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  exp_reg_5_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  exp_reg_5_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  exp_reg_6_0 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  exp_reg_6_1 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  exp_reg_7_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  exp_reg_7_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  exp_reg_8_0 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  exp_reg_8_1 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  new_frac_reg_0_0 = _RAND_28[23:0];
  _RAND_29 = {1{`RANDOM}};
  new_frac_reg_0_1 = _RAND_29[23:0];
  _RAND_30 = {1{`RANDOM}};
  new_frac_reg_1_0 = _RAND_30[23:0];
  _RAND_31 = {1{`RANDOM}};
  new_frac_reg_1_1 = _RAND_31[23:0];
  _RAND_32 = {2{`RANDOM}};
  multipplier_out_s_reg_0 = _RAND_32[47:0];
  _RAND_33 = {2{`RANDOM}};
  multipplier_out_s_reg_1 = _RAND_33[47:0];
  _RAND_34 = {2{`RANDOM}};
  multipplier_out_s_reg_2 = _RAND_34[47:0];
  _RAND_35 = {2{`RANDOM}};
  multipplier_out_s_reg_3 = _RAND_35[47:0];
  _RAND_36 = {2{`RANDOM}};
  multipplier_out_s_reg_4 = _RAND_36[47:0];
  _RAND_37 = {2{`RANDOM}};
  multipplier_out_s_reg_5 = _RAND_37[47:0];
  _RAND_38 = {1{`RANDOM}};
  subber_out_s_reg_0 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  complementN_out_reg_0 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  complementN_out_reg_1 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  complementN_out_reg_2 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  new_s_reg_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  new_s_reg_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  new_s_reg_2 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  new_s_reg_3 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  is_exp1_neg_reg_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  is_exp1_neg_reg_1 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  adderN_out_s_reg_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  adderN_out_c_reg_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  new_exp_reg_0 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  new_mant_reg_0 = _RAND_51[22:0];
  _RAND_52 = {1{`RANDOM}};
  reg_out_s = _RAND_52[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FP_reciprocal_newfpu(
  input         clock,
  input         reset,
  input         io_in_en,
  input  [31:0] io_in_a,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2077;
  reg [31:0] _RAND_2078;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [31:0] _RAND_2085;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [31:0] _RAND_2088;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [31:0] _RAND_2109;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [31:0] _RAND_2115;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2121;
  reg [31:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [31:0] _RAND_2124;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [31:0] _RAND_2163;
  reg [31:0] _RAND_2164;
  reg [31:0] _RAND_2165;
  reg [31:0] _RAND_2166;
  reg [31:0] _RAND_2167;
  reg [31:0] _RAND_2168;
  reg [31:0] _RAND_2169;
  reg [31:0] _RAND_2170;
  reg [31:0] _RAND_2171;
  reg [31:0] _RAND_2172;
  reg [31:0] _RAND_2173;
  reg [31:0] _RAND_2174;
  reg [31:0] _RAND_2175;
  reg [31:0] _RAND_2176;
  reg [31:0] _RAND_2177;
`endif // RANDOMIZE_REG_INIT
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_1_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_1_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_1_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_1_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_1_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_2_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_2_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_2_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_2_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_2_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_3_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_3_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_3_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_3_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_3_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_4_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_4_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_4_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_4_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_4_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_5_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_5_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_5_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_5_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_5_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_6_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_6_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_6_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_6_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_6_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_7_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_7_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_7_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_7_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_7_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_8_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_8_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_8_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_8_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_8_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_9_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_9_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_9_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_9_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_9_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_10_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_10_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_10_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_10_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_10_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_11_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_11_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_11_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_11_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_11_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_12_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_12_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_12_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_12_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_12_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_13_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_13_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_13_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_13_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_13_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_14_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_14_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_14_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_14_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_14_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_15_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_15_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_15_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_15_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_15_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_16_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_16_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_16_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_16_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_16_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_17_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_17_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_17_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_17_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_17_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_18_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_18_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_18_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_18_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_18_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_19_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_19_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_19_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_19_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_19_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_20_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_20_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_20_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_20_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_20_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_21_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_21_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_21_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_21_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_21_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_22_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_22_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_22_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_22_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_22_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_23_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_23_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_23_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_23_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_23_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_24_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_24_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_24_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_24_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_24_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_25_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_25_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_25_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_25_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_25_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_26_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_26_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_26_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_26_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_26_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_27_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_27_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_27_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_27_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_27_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_28_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_28_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_28_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_28_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_28_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_29_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_29_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_29_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_29_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_29_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_30_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_30_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_30_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_30_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_30_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_31_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_31_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_31_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_31_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_31_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_32_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_32_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_32_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_32_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_32_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_33_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_33_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_33_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_33_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_33_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_34_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_34_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_34_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_34_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_34_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_35_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_35_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_35_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_35_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_35_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_36_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_36_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_36_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_36_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_36_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_37_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_37_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_37_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_37_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_37_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_38_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_38_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_38_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_38_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_38_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_39_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_39_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_39_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_39_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_39_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_40_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_40_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_40_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_40_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_40_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_41_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_41_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_41_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_41_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_41_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_42_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_42_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_42_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_42_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_42_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_43_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_43_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_43_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_43_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_43_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_44_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_44_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_44_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_44_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_44_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_45_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_45_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_45_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_45_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_45_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_46_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_46_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_46_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_46_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_46_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_47_clock; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_47_reset; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_multiplier_10ccs_47_io_in_en; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_47_io_in_a; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_47_io_in_b; // @[FloatingPointDesigns.scala 2114:65]
  wire [31:0] FP_multiplier_10ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2114:65]
  wire  FP_subtractor_13ccs_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_1_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_1_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_1_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_1_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_1_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_2_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_2_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_2_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_2_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_2_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_3_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_3_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_3_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_3_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_3_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_4_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_4_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_4_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_4_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_4_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_5_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_5_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_5_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_5_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_5_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_6_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_6_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_6_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_6_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_6_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_7_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_7_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_7_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_7_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_7_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_8_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_8_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_8_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_8_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_8_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_9_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_9_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_9_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_9_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_9_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_10_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_10_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_10_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_10_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_10_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_11_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_11_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_11_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_11_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_11_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_12_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_12_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_12_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_12_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_12_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_13_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_13_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_13_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_13_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_13_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_14_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_14_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_14_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_14_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_14_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_15_clock; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_15_reset; // @[FloatingPointDesigns.scala 2115:50]
  wire  FP_subtractor_13ccs_15_io_in_en; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_15_io_in_a; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_15_io_in_b; // @[FloatingPointDesigns.scala 2115:50]
  wire [31:0] FP_subtractor_13ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2115:50]
  wire  multiplier4_clock; // @[FloatingPointDesigns.scala 2194:29]
  wire  multiplier4_reset; // @[FloatingPointDesigns.scala 2194:29]
  wire  multiplier4_io_in_en; // @[FloatingPointDesigns.scala 2194:29]
  wire [31:0] multiplier4_io_in_a; // @[FloatingPointDesigns.scala 2194:29]
  wire [31:0] multiplier4_io_in_b; // @[FloatingPointDesigns.scala 2194:29]
  wire [31:0] multiplier4_io_out_s; // @[FloatingPointDesigns.scala 2194:29]
  wire  FP_multiplier_10ccs_48_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_48_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_48_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_48_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_48_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_49_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_49_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_49_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_49_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_49_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_50_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_50_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_50_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_50_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_50_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_51_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_51_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_51_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_51_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_51_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_52_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_52_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_52_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_52_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_52_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_53_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_53_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_53_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_53_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_53_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_54_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_54_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_54_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_54_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_54_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_55_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_55_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_55_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_55_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_55_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_56_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_56_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_56_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_56_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_56_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_57_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_57_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_57_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_57_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_57_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_58_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_58_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_58_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_58_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_58_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_59_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_59_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_59_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_59_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_59_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_60_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_60_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_60_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_60_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_60_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_61_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_61_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_61_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_61_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_61_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_62_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_62_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_62_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_62_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_62_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_63_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_63_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_63_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_63_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_63_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_64_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_64_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_64_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_64_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_64_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_64_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_65_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_65_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_65_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_65_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_65_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_65_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_66_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_66_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_66_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_66_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_66_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_66_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_67_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_67_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_67_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_67_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_67_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_67_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_68_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_68_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_68_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_68_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_68_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_68_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_69_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_69_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_69_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_69_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_69_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_69_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_70_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_70_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_70_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_70_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_70_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_70_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_71_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_71_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_71_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_71_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_71_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_71_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_72_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_72_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_72_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_72_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_72_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_72_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_73_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_73_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_73_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_73_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_73_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_73_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_74_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_74_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_74_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_74_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_74_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_74_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_75_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_75_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_75_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_75_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_75_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_75_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_76_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_76_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_76_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_76_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_76_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_76_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_77_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_77_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_77_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_77_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_77_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_77_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_78_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_78_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_78_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_78_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_78_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_78_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_79_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_79_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_79_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_79_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_79_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_79_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_80_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_80_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_80_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_80_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_80_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_80_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_81_clock; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_81_reset; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_multiplier_10ccs_81_io_in_en; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_81_io_in_a; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_81_io_in_b; // @[FloatingPointDesigns.scala 2206:69]
  wire [31:0] FP_multiplier_10ccs_81_io_out_s; // @[FloatingPointDesigns.scala 2206:69]
  wire  FP_subtractor_13ccs_16_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_16_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_16_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_16_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_16_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_17_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_17_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_17_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_17_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_17_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_18_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_18_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_18_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_18_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_18_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_19_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_19_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_19_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_19_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_19_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_20_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_20_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_20_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_20_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_20_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_21_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_21_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_21_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_21_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_21_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_22_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_22_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_22_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_22_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_22_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_23_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_23_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_23_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_23_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_23_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_24_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_24_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_24_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_24_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_24_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_25_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_25_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_25_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_25_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_25_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_26_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_26_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_26_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_26_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_26_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_27_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_27_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_27_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_27_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_27_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_28_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_28_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_28_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_28_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_28_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_29_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_29_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_29_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_29_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_29_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_30_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_30_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_30_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_30_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_30_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_31_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_31_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_31_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_31_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_31_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_32_clock; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_32_reset; // @[FloatingPointDesigns.scala 2207:54]
  wire  FP_subtractor_13ccs_32_io_in_en; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_32_io_in_a; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_32_io_in_b; // @[FloatingPointDesigns.scala 2207:54]
  wire [31:0] FP_subtractor_13ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2207:54]
  wire [30:0] _number_T_1 = {{1'd0}, io_in_a[30:1]}; // @[FloatingPointDesigns.scala 2099:36]
  wire [30:0] _GEN_0 = io_in_a[30:0] > 31'h7ef477d4 ? 31'h3f7a3bea : _number_T_1; // @[FloatingPointDesigns.scala 2096:46 2097:14 2099:14]
  wire [31:0] number = {{1'd0}, _GEN_0}; // @[FloatingPointDesigns.scala 2091:22]
  wire [31:0] result = 32'h5f3759df - number; // @[FloatingPointDesigns.scala 2106:25]
  reg [31:0] x_n_0; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_1; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_2; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_4; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_5; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_6; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_8; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_9; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_10; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_12; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_13; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_14; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_16; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_17; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_18; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_20; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_21; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_22; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_24; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_25; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_26; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_28; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_29; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_30; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_32; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_33; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_34; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_36; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_37; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_38; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_40; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_41; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_42; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_44; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_45; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_46; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_48; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_49; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_50; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_52; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_53; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_54; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_56; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_57; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_58; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_60; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_61; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] x_n_62; // @[FloatingPointDesigns.scala 2108:22]
  reg [31:0] a_2_0; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_1; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_2; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_3; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_4; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_5; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_6; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_7; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_8; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_9; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_10; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_11; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_12; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_13; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_14; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_15; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_16; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_17; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_18; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_19; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_20; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_21; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_22; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_23; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_24; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_25; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_26; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_27; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_28; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_29; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_30; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_31; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_32; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_33; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_34; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_35; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_36; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_37; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_38; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_39; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_40; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_41; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_42; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_43; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_44; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_45; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_46; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_47; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_48; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_49; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_50; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_51; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_52; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_53; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_54; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_55; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_56; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_57; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_58; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_59; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_60; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_61; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_62; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] a_2_63; // @[FloatingPointDesigns.scala 2109:22]
  reg [31:0] stage1_regs_0_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_0_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_1_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_2_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_3_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_4_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_5_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_6_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_7_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_8_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_9_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_10_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_11_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_12_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_13_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_14_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_0_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_0_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_0_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_0_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_0_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_0_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_0_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_0_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_0_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_1_0; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_1_1; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_1_2; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_1_3; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_1_4; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_1_5; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_1_6; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_1_7; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage1_regs_15_1_8; // @[FloatingPointDesigns.scala 2110:30]
  reg [31:0] stage2_regs_0_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_0_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_1_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_2_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_3_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_4_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_5_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_6_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_7_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_8_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_9_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_10_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_11_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_12_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_13_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_14_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_0_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_0_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_0_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_0_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_0_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_0_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_0_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_0_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_0_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_1_0; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_1_1; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_1_2; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_1_3; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_1_4; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_1_5; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_1_6; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_1_7; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage2_regs_15_1_8; // @[FloatingPointDesigns.scala 2111:30]
  reg [31:0] stage3_regs_0_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_0_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_1_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_2_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_3_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_4_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_5_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_6_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_7_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_8_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_9_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_10_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_11_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_12_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_13_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_14_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_0_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_0_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_0_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_0_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_0_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_0_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_0_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_0_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_0_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_0_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_0_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_0_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_1_0; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_1_1; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_1_2; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_1_3; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_1_4; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_1_5; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_1_6; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_1_7; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_1_8; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_1_9; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_1_10; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage3_regs_15_1_11; // @[FloatingPointDesigns.scala 2112:30]
  reg [31:0] stage4_regs_0_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_0_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_0_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_0_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_0_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_0_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_0_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_0_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_0_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_1_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_1_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_1_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_1_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_1_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_1_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_1_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_1_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_1_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_2_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_2_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_2_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_2_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_2_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_2_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_2_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_2_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_2_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_3_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_3_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_3_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_3_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_3_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_3_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_3_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_3_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_3_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_4_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_4_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_4_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_4_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_4_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_4_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_4_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_4_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_4_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_5_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_5_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_5_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_5_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_5_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_5_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_5_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_5_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_5_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_6_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_6_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_6_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_6_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_6_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_6_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_6_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_6_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_6_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_7_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_7_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_7_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_7_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_7_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_7_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_7_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_7_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_7_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_8_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_8_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_8_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_8_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_8_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_8_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_8_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_8_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_8_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_9_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_9_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_9_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_9_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_9_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_9_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_9_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_9_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_9_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_10_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_10_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_10_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_10_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_10_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_10_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_10_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_10_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_10_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_11_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_11_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_11_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_11_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_11_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_11_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_11_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_11_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_11_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_12_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_12_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_12_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_12_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_12_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_12_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_12_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_12_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_12_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_13_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_13_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_13_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_13_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_13_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_13_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_13_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_13_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_13_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_14_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_14_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_14_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_14_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_14_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_14_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_14_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_14_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_14_1_8; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_15_1_0; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_15_1_1; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_15_1_2; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_15_1_3; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_15_1_4; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_15_1_5; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_15_1_6; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_15_1_7; // @[FloatingPointDesigns.scala 2113:30]
  reg [31:0] stage4_regs_15_1_8; // @[FloatingPointDesigns.scala 2113:30]
  wire [7:0] _a_2_0_T_3 = io_in_a[30:23] - 8'h1; // @[FloatingPointDesigns.scala 2139:75]
  wire [31:0] _a_2_0_T_6 = {io_in_a[31],_a_2_0_T_3,io_in_a[22:0]}; // @[FloatingPointDesigns.scala 2139:82]
  reg [31:0] a_2_isr_to_r; // @[FloatingPointDesigns.scala 2184:31]
  reg [31:0] transition_regs_0; // @[FloatingPointDesigns.scala 2185:34]
  reg [31:0] transition_regs_1; // @[FloatingPointDesigns.scala 2185:34]
  reg [31:0] transition_regs_2; // @[FloatingPointDesigns.scala 2185:34]
  reg [31:0] transition_regs_3; // @[FloatingPointDesigns.scala 2185:34]
  reg [31:0] transition_regs_4; // @[FloatingPointDesigns.scala 2185:34]
  reg [31:0] transition_regs_5; // @[FloatingPointDesigns.scala 2185:34]
  reg [31:0] transition_regs_6; // @[FloatingPointDesigns.scala 2185:34]
  reg [31:0] transition_regs_7; // @[FloatingPointDesigns.scala 2185:34]
  reg [31:0] transition_regs_8; // @[FloatingPointDesigns.scala 2185:34]
  wire [7:0] _a_2_isr_to_r_T_3 = stage4_regs_15_1_8[30:23] + 8'h1; // @[FloatingPointDesigns.scala 2187:115]
  wire [31:0] _a_2_isr_to_r_T_6 = {stage4_regs_15_1_8[31],_a_2_isr_to_r_T_3,stage4_regs_15_1_8[22:0]}; // @[FloatingPointDesigns.scala 2187:122]
  reg [31:0] x_n_r_0; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_1; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_3; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_4; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_6; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_7; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_9; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_10; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_12; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_13; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_15; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_16; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_18; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_19; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_21; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_22; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_24; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_25; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_27; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_28; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_30; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_31; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_33; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_34; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_36; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_37; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_39; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_40; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_42; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_43; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_45; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_46; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_48; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] x_n_r_49; // @[FloatingPointDesigns.scala 2201:24]
  reg [31:0] a_2_r_0; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_1; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_2; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_3; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_4; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_5; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_6; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_7; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_8; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_9; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_10; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_11; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_12; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_13; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_14; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_15; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_16; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_17; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_18; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_19; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_20; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_21; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_22; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_23; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_24; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_25; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_26; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_27; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_28; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_29; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_30; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_31; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_32; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_33; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_34; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_35; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_36; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_37; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_38; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_39; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_40; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_41; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_42; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_43; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_44; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_45; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_46; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_47; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_48; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_49; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] a_2_r_50; // @[FloatingPointDesigns.scala 2202:24]
  reg [31:0] stage1_regs_r_0_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_0_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_1_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_2_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_3_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_4_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_5_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_6_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_7_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_8_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_9_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_10_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_11_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_12_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_13_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_14_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_15_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_0_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_0_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_0_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_0_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_0_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_0_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_0_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_0_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_0_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_1_0; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_1_1; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_1_2; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_1_3; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_1_4; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_1_5; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_1_6; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_1_7; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage1_regs_r_16_1_8; // @[FloatingPointDesigns.scala 2203:32]
  reg [31:0] stage2_regs_r_0_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_0_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_1_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_2_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_3_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_4_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_5_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_6_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_7_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_8_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_9_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_10_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_11_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_12_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_13_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_14_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_15_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_0_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_0_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_0_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_0_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_0_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_0_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_0_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_0_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_0_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_0_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_0_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_0_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_1_0; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_1_1; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_1_2; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_1_3; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_1_4; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_1_5; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_1_6; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_1_7; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_1_8; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_1_9; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_1_10; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage2_regs_r_16_1_11; // @[FloatingPointDesigns.scala 2204:32]
  reg [31:0] stage3_regs_r_0_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_0_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_0_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_0_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_0_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_0_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_0_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_0_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_0_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_1_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_1_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_1_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_1_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_1_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_1_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_1_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_1_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_1_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_2_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_2_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_2_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_2_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_2_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_2_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_2_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_2_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_2_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_3_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_3_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_3_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_3_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_3_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_3_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_3_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_3_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_3_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_4_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_4_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_4_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_4_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_4_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_4_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_4_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_4_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_4_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_5_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_5_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_5_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_5_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_5_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_5_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_5_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_5_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_5_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_6_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_6_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_6_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_6_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_6_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_6_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_6_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_6_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_6_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_7_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_7_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_7_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_7_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_7_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_7_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_7_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_7_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_7_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_8_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_8_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_8_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_8_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_8_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_8_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_8_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_8_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_8_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_9_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_9_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_9_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_9_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_9_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_9_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_9_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_9_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_9_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_10_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_10_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_10_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_10_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_10_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_10_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_10_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_10_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_10_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_11_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_11_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_11_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_11_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_11_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_11_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_11_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_11_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_11_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_12_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_12_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_12_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_12_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_12_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_12_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_12_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_12_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_12_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_13_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_13_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_13_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_13_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_13_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_13_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_13_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_13_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_13_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_14_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_14_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_14_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_14_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_14_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_14_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_14_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_14_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_14_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_15_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_15_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_15_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_15_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_15_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_15_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_15_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_15_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_15_1_8; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_16_1_0; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_16_1_1; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_16_1_2; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_16_1_3; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_16_1_4; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_16_1_5; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_16_1_6; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_16_1_7; // @[FloatingPointDesigns.scala 2205:32]
  reg [31:0] stage3_regs_r_16_1_8; // @[FloatingPointDesigns.scala 2205:32]
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_en(FP_multiplier_10ccs_io_in_en),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_1 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_1_clock),
    .reset(FP_multiplier_10ccs_1_reset),
    .io_in_en(FP_multiplier_10ccs_1_io_in_en),
    .io_in_a(FP_multiplier_10ccs_1_io_in_a),
    .io_in_b(FP_multiplier_10ccs_1_io_in_b),
    .io_out_s(FP_multiplier_10ccs_1_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_2 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_2_clock),
    .reset(FP_multiplier_10ccs_2_reset),
    .io_in_en(FP_multiplier_10ccs_2_io_in_en),
    .io_in_a(FP_multiplier_10ccs_2_io_in_a),
    .io_in_b(FP_multiplier_10ccs_2_io_in_b),
    .io_out_s(FP_multiplier_10ccs_2_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_3 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_3_clock),
    .reset(FP_multiplier_10ccs_3_reset),
    .io_in_en(FP_multiplier_10ccs_3_io_in_en),
    .io_in_a(FP_multiplier_10ccs_3_io_in_a),
    .io_in_b(FP_multiplier_10ccs_3_io_in_b),
    .io_out_s(FP_multiplier_10ccs_3_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_4 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_4_clock),
    .reset(FP_multiplier_10ccs_4_reset),
    .io_in_en(FP_multiplier_10ccs_4_io_in_en),
    .io_in_a(FP_multiplier_10ccs_4_io_in_a),
    .io_in_b(FP_multiplier_10ccs_4_io_in_b),
    .io_out_s(FP_multiplier_10ccs_4_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_5 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_5_clock),
    .reset(FP_multiplier_10ccs_5_reset),
    .io_in_en(FP_multiplier_10ccs_5_io_in_en),
    .io_in_a(FP_multiplier_10ccs_5_io_in_a),
    .io_in_b(FP_multiplier_10ccs_5_io_in_b),
    .io_out_s(FP_multiplier_10ccs_5_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_6 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_6_clock),
    .reset(FP_multiplier_10ccs_6_reset),
    .io_in_en(FP_multiplier_10ccs_6_io_in_en),
    .io_in_a(FP_multiplier_10ccs_6_io_in_a),
    .io_in_b(FP_multiplier_10ccs_6_io_in_b),
    .io_out_s(FP_multiplier_10ccs_6_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_7 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_7_clock),
    .reset(FP_multiplier_10ccs_7_reset),
    .io_in_en(FP_multiplier_10ccs_7_io_in_en),
    .io_in_a(FP_multiplier_10ccs_7_io_in_a),
    .io_in_b(FP_multiplier_10ccs_7_io_in_b),
    .io_out_s(FP_multiplier_10ccs_7_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_8 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_8_clock),
    .reset(FP_multiplier_10ccs_8_reset),
    .io_in_en(FP_multiplier_10ccs_8_io_in_en),
    .io_in_a(FP_multiplier_10ccs_8_io_in_a),
    .io_in_b(FP_multiplier_10ccs_8_io_in_b),
    .io_out_s(FP_multiplier_10ccs_8_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_9 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_9_clock),
    .reset(FP_multiplier_10ccs_9_reset),
    .io_in_en(FP_multiplier_10ccs_9_io_in_en),
    .io_in_a(FP_multiplier_10ccs_9_io_in_a),
    .io_in_b(FP_multiplier_10ccs_9_io_in_b),
    .io_out_s(FP_multiplier_10ccs_9_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_10 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_10_clock),
    .reset(FP_multiplier_10ccs_10_reset),
    .io_in_en(FP_multiplier_10ccs_10_io_in_en),
    .io_in_a(FP_multiplier_10ccs_10_io_in_a),
    .io_in_b(FP_multiplier_10ccs_10_io_in_b),
    .io_out_s(FP_multiplier_10ccs_10_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_11 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_11_clock),
    .reset(FP_multiplier_10ccs_11_reset),
    .io_in_en(FP_multiplier_10ccs_11_io_in_en),
    .io_in_a(FP_multiplier_10ccs_11_io_in_a),
    .io_in_b(FP_multiplier_10ccs_11_io_in_b),
    .io_out_s(FP_multiplier_10ccs_11_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_12 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_12_clock),
    .reset(FP_multiplier_10ccs_12_reset),
    .io_in_en(FP_multiplier_10ccs_12_io_in_en),
    .io_in_a(FP_multiplier_10ccs_12_io_in_a),
    .io_in_b(FP_multiplier_10ccs_12_io_in_b),
    .io_out_s(FP_multiplier_10ccs_12_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_13 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_13_clock),
    .reset(FP_multiplier_10ccs_13_reset),
    .io_in_en(FP_multiplier_10ccs_13_io_in_en),
    .io_in_a(FP_multiplier_10ccs_13_io_in_a),
    .io_in_b(FP_multiplier_10ccs_13_io_in_b),
    .io_out_s(FP_multiplier_10ccs_13_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_14 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_14_clock),
    .reset(FP_multiplier_10ccs_14_reset),
    .io_in_en(FP_multiplier_10ccs_14_io_in_en),
    .io_in_a(FP_multiplier_10ccs_14_io_in_a),
    .io_in_b(FP_multiplier_10ccs_14_io_in_b),
    .io_out_s(FP_multiplier_10ccs_14_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_15 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_15_clock),
    .reset(FP_multiplier_10ccs_15_reset),
    .io_in_en(FP_multiplier_10ccs_15_io_in_en),
    .io_in_a(FP_multiplier_10ccs_15_io_in_a),
    .io_in_b(FP_multiplier_10ccs_15_io_in_b),
    .io_out_s(FP_multiplier_10ccs_15_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_16 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_16_clock),
    .reset(FP_multiplier_10ccs_16_reset),
    .io_in_en(FP_multiplier_10ccs_16_io_in_en),
    .io_in_a(FP_multiplier_10ccs_16_io_in_a),
    .io_in_b(FP_multiplier_10ccs_16_io_in_b),
    .io_out_s(FP_multiplier_10ccs_16_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_17 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_17_clock),
    .reset(FP_multiplier_10ccs_17_reset),
    .io_in_en(FP_multiplier_10ccs_17_io_in_en),
    .io_in_a(FP_multiplier_10ccs_17_io_in_a),
    .io_in_b(FP_multiplier_10ccs_17_io_in_b),
    .io_out_s(FP_multiplier_10ccs_17_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_18 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_18_clock),
    .reset(FP_multiplier_10ccs_18_reset),
    .io_in_en(FP_multiplier_10ccs_18_io_in_en),
    .io_in_a(FP_multiplier_10ccs_18_io_in_a),
    .io_in_b(FP_multiplier_10ccs_18_io_in_b),
    .io_out_s(FP_multiplier_10ccs_18_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_19 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_19_clock),
    .reset(FP_multiplier_10ccs_19_reset),
    .io_in_en(FP_multiplier_10ccs_19_io_in_en),
    .io_in_a(FP_multiplier_10ccs_19_io_in_a),
    .io_in_b(FP_multiplier_10ccs_19_io_in_b),
    .io_out_s(FP_multiplier_10ccs_19_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_20 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_20_clock),
    .reset(FP_multiplier_10ccs_20_reset),
    .io_in_en(FP_multiplier_10ccs_20_io_in_en),
    .io_in_a(FP_multiplier_10ccs_20_io_in_a),
    .io_in_b(FP_multiplier_10ccs_20_io_in_b),
    .io_out_s(FP_multiplier_10ccs_20_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_21 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_21_clock),
    .reset(FP_multiplier_10ccs_21_reset),
    .io_in_en(FP_multiplier_10ccs_21_io_in_en),
    .io_in_a(FP_multiplier_10ccs_21_io_in_a),
    .io_in_b(FP_multiplier_10ccs_21_io_in_b),
    .io_out_s(FP_multiplier_10ccs_21_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_22 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_22_clock),
    .reset(FP_multiplier_10ccs_22_reset),
    .io_in_en(FP_multiplier_10ccs_22_io_in_en),
    .io_in_a(FP_multiplier_10ccs_22_io_in_a),
    .io_in_b(FP_multiplier_10ccs_22_io_in_b),
    .io_out_s(FP_multiplier_10ccs_22_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_23 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_23_clock),
    .reset(FP_multiplier_10ccs_23_reset),
    .io_in_en(FP_multiplier_10ccs_23_io_in_en),
    .io_in_a(FP_multiplier_10ccs_23_io_in_a),
    .io_in_b(FP_multiplier_10ccs_23_io_in_b),
    .io_out_s(FP_multiplier_10ccs_23_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_24 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_24_clock),
    .reset(FP_multiplier_10ccs_24_reset),
    .io_in_en(FP_multiplier_10ccs_24_io_in_en),
    .io_in_a(FP_multiplier_10ccs_24_io_in_a),
    .io_in_b(FP_multiplier_10ccs_24_io_in_b),
    .io_out_s(FP_multiplier_10ccs_24_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_25 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_25_clock),
    .reset(FP_multiplier_10ccs_25_reset),
    .io_in_en(FP_multiplier_10ccs_25_io_in_en),
    .io_in_a(FP_multiplier_10ccs_25_io_in_a),
    .io_in_b(FP_multiplier_10ccs_25_io_in_b),
    .io_out_s(FP_multiplier_10ccs_25_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_26 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_26_clock),
    .reset(FP_multiplier_10ccs_26_reset),
    .io_in_en(FP_multiplier_10ccs_26_io_in_en),
    .io_in_a(FP_multiplier_10ccs_26_io_in_a),
    .io_in_b(FP_multiplier_10ccs_26_io_in_b),
    .io_out_s(FP_multiplier_10ccs_26_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_27 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_27_clock),
    .reset(FP_multiplier_10ccs_27_reset),
    .io_in_en(FP_multiplier_10ccs_27_io_in_en),
    .io_in_a(FP_multiplier_10ccs_27_io_in_a),
    .io_in_b(FP_multiplier_10ccs_27_io_in_b),
    .io_out_s(FP_multiplier_10ccs_27_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_28 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_28_clock),
    .reset(FP_multiplier_10ccs_28_reset),
    .io_in_en(FP_multiplier_10ccs_28_io_in_en),
    .io_in_a(FP_multiplier_10ccs_28_io_in_a),
    .io_in_b(FP_multiplier_10ccs_28_io_in_b),
    .io_out_s(FP_multiplier_10ccs_28_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_29 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_29_clock),
    .reset(FP_multiplier_10ccs_29_reset),
    .io_in_en(FP_multiplier_10ccs_29_io_in_en),
    .io_in_a(FP_multiplier_10ccs_29_io_in_a),
    .io_in_b(FP_multiplier_10ccs_29_io_in_b),
    .io_out_s(FP_multiplier_10ccs_29_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_30 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_30_clock),
    .reset(FP_multiplier_10ccs_30_reset),
    .io_in_en(FP_multiplier_10ccs_30_io_in_en),
    .io_in_a(FP_multiplier_10ccs_30_io_in_a),
    .io_in_b(FP_multiplier_10ccs_30_io_in_b),
    .io_out_s(FP_multiplier_10ccs_30_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_31 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_31_clock),
    .reset(FP_multiplier_10ccs_31_reset),
    .io_in_en(FP_multiplier_10ccs_31_io_in_en),
    .io_in_a(FP_multiplier_10ccs_31_io_in_a),
    .io_in_b(FP_multiplier_10ccs_31_io_in_b),
    .io_out_s(FP_multiplier_10ccs_31_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_32 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_32_clock),
    .reset(FP_multiplier_10ccs_32_reset),
    .io_in_en(FP_multiplier_10ccs_32_io_in_en),
    .io_in_a(FP_multiplier_10ccs_32_io_in_a),
    .io_in_b(FP_multiplier_10ccs_32_io_in_b),
    .io_out_s(FP_multiplier_10ccs_32_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_33 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_33_clock),
    .reset(FP_multiplier_10ccs_33_reset),
    .io_in_en(FP_multiplier_10ccs_33_io_in_en),
    .io_in_a(FP_multiplier_10ccs_33_io_in_a),
    .io_in_b(FP_multiplier_10ccs_33_io_in_b),
    .io_out_s(FP_multiplier_10ccs_33_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_34 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_34_clock),
    .reset(FP_multiplier_10ccs_34_reset),
    .io_in_en(FP_multiplier_10ccs_34_io_in_en),
    .io_in_a(FP_multiplier_10ccs_34_io_in_a),
    .io_in_b(FP_multiplier_10ccs_34_io_in_b),
    .io_out_s(FP_multiplier_10ccs_34_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_35 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_35_clock),
    .reset(FP_multiplier_10ccs_35_reset),
    .io_in_en(FP_multiplier_10ccs_35_io_in_en),
    .io_in_a(FP_multiplier_10ccs_35_io_in_a),
    .io_in_b(FP_multiplier_10ccs_35_io_in_b),
    .io_out_s(FP_multiplier_10ccs_35_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_36 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_36_clock),
    .reset(FP_multiplier_10ccs_36_reset),
    .io_in_en(FP_multiplier_10ccs_36_io_in_en),
    .io_in_a(FP_multiplier_10ccs_36_io_in_a),
    .io_in_b(FP_multiplier_10ccs_36_io_in_b),
    .io_out_s(FP_multiplier_10ccs_36_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_37 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_37_clock),
    .reset(FP_multiplier_10ccs_37_reset),
    .io_in_en(FP_multiplier_10ccs_37_io_in_en),
    .io_in_a(FP_multiplier_10ccs_37_io_in_a),
    .io_in_b(FP_multiplier_10ccs_37_io_in_b),
    .io_out_s(FP_multiplier_10ccs_37_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_38 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_38_clock),
    .reset(FP_multiplier_10ccs_38_reset),
    .io_in_en(FP_multiplier_10ccs_38_io_in_en),
    .io_in_a(FP_multiplier_10ccs_38_io_in_a),
    .io_in_b(FP_multiplier_10ccs_38_io_in_b),
    .io_out_s(FP_multiplier_10ccs_38_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_39 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_39_clock),
    .reset(FP_multiplier_10ccs_39_reset),
    .io_in_en(FP_multiplier_10ccs_39_io_in_en),
    .io_in_a(FP_multiplier_10ccs_39_io_in_a),
    .io_in_b(FP_multiplier_10ccs_39_io_in_b),
    .io_out_s(FP_multiplier_10ccs_39_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_40 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_40_clock),
    .reset(FP_multiplier_10ccs_40_reset),
    .io_in_en(FP_multiplier_10ccs_40_io_in_en),
    .io_in_a(FP_multiplier_10ccs_40_io_in_a),
    .io_in_b(FP_multiplier_10ccs_40_io_in_b),
    .io_out_s(FP_multiplier_10ccs_40_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_41 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_41_clock),
    .reset(FP_multiplier_10ccs_41_reset),
    .io_in_en(FP_multiplier_10ccs_41_io_in_en),
    .io_in_a(FP_multiplier_10ccs_41_io_in_a),
    .io_in_b(FP_multiplier_10ccs_41_io_in_b),
    .io_out_s(FP_multiplier_10ccs_41_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_42 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_42_clock),
    .reset(FP_multiplier_10ccs_42_reset),
    .io_in_en(FP_multiplier_10ccs_42_io_in_en),
    .io_in_a(FP_multiplier_10ccs_42_io_in_a),
    .io_in_b(FP_multiplier_10ccs_42_io_in_b),
    .io_out_s(FP_multiplier_10ccs_42_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_43 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_43_clock),
    .reset(FP_multiplier_10ccs_43_reset),
    .io_in_en(FP_multiplier_10ccs_43_io_in_en),
    .io_in_a(FP_multiplier_10ccs_43_io_in_a),
    .io_in_b(FP_multiplier_10ccs_43_io_in_b),
    .io_out_s(FP_multiplier_10ccs_43_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_44 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_44_clock),
    .reset(FP_multiplier_10ccs_44_reset),
    .io_in_en(FP_multiplier_10ccs_44_io_in_en),
    .io_in_a(FP_multiplier_10ccs_44_io_in_a),
    .io_in_b(FP_multiplier_10ccs_44_io_in_b),
    .io_out_s(FP_multiplier_10ccs_44_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_45 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_45_clock),
    .reset(FP_multiplier_10ccs_45_reset),
    .io_in_en(FP_multiplier_10ccs_45_io_in_en),
    .io_in_a(FP_multiplier_10ccs_45_io_in_a),
    .io_in_b(FP_multiplier_10ccs_45_io_in_b),
    .io_out_s(FP_multiplier_10ccs_45_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_46 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_46_clock),
    .reset(FP_multiplier_10ccs_46_reset),
    .io_in_en(FP_multiplier_10ccs_46_io_in_en),
    .io_in_a(FP_multiplier_10ccs_46_io_in_a),
    .io_in_b(FP_multiplier_10ccs_46_io_in_b),
    .io_out_s(FP_multiplier_10ccs_46_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_47 ( // @[FloatingPointDesigns.scala 2114:65]
    .clock(FP_multiplier_10ccs_47_clock),
    .reset(FP_multiplier_10ccs_47_reset),
    .io_in_en(FP_multiplier_10ccs_47_io_in_en),
    .io_in_a(FP_multiplier_10ccs_47_io_in_a),
    .io_in_b(FP_multiplier_10ccs_47_io_in_b),
    .io_out_s(FP_multiplier_10ccs_47_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_clock),
    .reset(FP_subtractor_13ccs_reset),
    .io_in_en(FP_subtractor_13ccs_io_in_en),
    .io_in_a(FP_subtractor_13ccs_io_in_a),
    .io_in_b(FP_subtractor_13ccs_io_in_b),
    .io_out_s(FP_subtractor_13ccs_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_1 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_1_clock),
    .reset(FP_subtractor_13ccs_1_reset),
    .io_in_en(FP_subtractor_13ccs_1_io_in_en),
    .io_in_a(FP_subtractor_13ccs_1_io_in_a),
    .io_in_b(FP_subtractor_13ccs_1_io_in_b),
    .io_out_s(FP_subtractor_13ccs_1_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_2 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_2_clock),
    .reset(FP_subtractor_13ccs_2_reset),
    .io_in_en(FP_subtractor_13ccs_2_io_in_en),
    .io_in_a(FP_subtractor_13ccs_2_io_in_a),
    .io_in_b(FP_subtractor_13ccs_2_io_in_b),
    .io_out_s(FP_subtractor_13ccs_2_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_3 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_3_clock),
    .reset(FP_subtractor_13ccs_3_reset),
    .io_in_en(FP_subtractor_13ccs_3_io_in_en),
    .io_in_a(FP_subtractor_13ccs_3_io_in_a),
    .io_in_b(FP_subtractor_13ccs_3_io_in_b),
    .io_out_s(FP_subtractor_13ccs_3_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_4 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_4_clock),
    .reset(FP_subtractor_13ccs_4_reset),
    .io_in_en(FP_subtractor_13ccs_4_io_in_en),
    .io_in_a(FP_subtractor_13ccs_4_io_in_a),
    .io_in_b(FP_subtractor_13ccs_4_io_in_b),
    .io_out_s(FP_subtractor_13ccs_4_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_5 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_5_clock),
    .reset(FP_subtractor_13ccs_5_reset),
    .io_in_en(FP_subtractor_13ccs_5_io_in_en),
    .io_in_a(FP_subtractor_13ccs_5_io_in_a),
    .io_in_b(FP_subtractor_13ccs_5_io_in_b),
    .io_out_s(FP_subtractor_13ccs_5_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_6 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_6_clock),
    .reset(FP_subtractor_13ccs_6_reset),
    .io_in_en(FP_subtractor_13ccs_6_io_in_en),
    .io_in_a(FP_subtractor_13ccs_6_io_in_a),
    .io_in_b(FP_subtractor_13ccs_6_io_in_b),
    .io_out_s(FP_subtractor_13ccs_6_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_7 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_7_clock),
    .reset(FP_subtractor_13ccs_7_reset),
    .io_in_en(FP_subtractor_13ccs_7_io_in_en),
    .io_in_a(FP_subtractor_13ccs_7_io_in_a),
    .io_in_b(FP_subtractor_13ccs_7_io_in_b),
    .io_out_s(FP_subtractor_13ccs_7_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_8 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_8_clock),
    .reset(FP_subtractor_13ccs_8_reset),
    .io_in_en(FP_subtractor_13ccs_8_io_in_en),
    .io_in_a(FP_subtractor_13ccs_8_io_in_a),
    .io_in_b(FP_subtractor_13ccs_8_io_in_b),
    .io_out_s(FP_subtractor_13ccs_8_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_9 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_9_clock),
    .reset(FP_subtractor_13ccs_9_reset),
    .io_in_en(FP_subtractor_13ccs_9_io_in_en),
    .io_in_a(FP_subtractor_13ccs_9_io_in_a),
    .io_in_b(FP_subtractor_13ccs_9_io_in_b),
    .io_out_s(FP_subtractor_13ccs_9_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_10 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_10_clock),
    .reset(FP_subtractor_13ccs_10_reset),
    .io_in_en(FP_subtractor_13ccs_10_io_in_en),
    .io_in_a(FP_subtractor_13ccs_10_io_in_a),
    .io_in_b(FP_subtractor_13ccs_10_io_in_b),
    .io_out_s(FP_subtractor_13ccs_10_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_11 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_11_clock),
    .reset(FP_subtractor_13ccs_11_reset),
    .io_in_en(FP_subtractor_13ccs_11_io_in_en),
    .io_in_a(FP_subtractor_13ccs_11_io_in_a),
    .io_in_b(FP_subtractor_13ccs_11_io_in_b),
    .io_out_s(FP_subtractor_13ccs_11_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_12 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_12_clock),
    .reset(FP_subtractor_13ccs_12_reset),
    .io_in_en(FP_subtractor_13ccs_12_io_in_en),
    .io_in_a(FP_subtractor_13ccs_12_io_in_a),
    .io_in_b(FP_subtractor_13ccs_12_io_in_b),
    .io_out_s(FP_subtractor_13ccs_12_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_13 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_13_clock),
    .reset(FP_subtractor_13ccs_13_reset),
    .io_in_en(FP_subtractor_13ccs_13_io_in_en),
    .io_in_a(FP_subtractor_13ccs_13_io_in_a),
    .io_in_b(FP_subtractor_13ccs_13_io_in_b),
    .io_out_s(FP_subtractor_13ccs_13_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_14 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_14_clock),
    .reset(FP_subtractor_13ccs_14_reset),
    .io_in_en(FP_subtractor_13ccs_14_io_in_en),
    .io_in_a(FP_subtractor_13ccs_14_io_in_a),
    .io_in_b(FP_subtractor_13ccs_14_io_in_b),
    .io_out_s(FP_subtractor_13ccs_14_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_15 ( // @[FloatingPointDesigns.scala 2115:50]
    .clock(FP_subtractor_13ccs_15_clock),
    .reset(FP_subtractor_13ccs_15_reset),
    .io_in_en(FP_subtractor_13ccs_15_io_in_en),
    .io_in_a(FP_subtractor_13ccs_15_io_in_a),
    .io_in_b(FP_subtractor_13ccs_15_io_in_b),
    .io_out_s(FP_subtractor_13ccs_15_io_out_s)
  );
  FP_multiplier_10ccs multiplier4 ( // @[FloatingPointDesigns.scala 2194:29]
    .clock(multiplier4_clock),
    .reset(multiplier4_reset),
    .io_in_en(multiplier4_io_in_en),
    .io_in_a(multiplier4_io_in_a),
    .io_in_b(multiplier4_io_in_b),
    .io_out_s(multiplier4_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_48 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_48_clock),
    .reset(FP_multiplier_10ccs_48_reset),
    .io_in_en(FP_multiplier_10ccs_48_io_in_en),
    .io_in_a(FP_multiplier_10ccs_48_io_in_a),
    .io_in_b(FP_multiplier_10ccs_48_io_in_b),
    .io_out_s(FP_multiplier_10ccs_48_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_49 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_49_clock),
    .reset(FP_multiplier_10ccs_49_reset),
    .io_in_en(FP_multiplier_10ccs_49_io_in_en),
    .io_in_a(FP_multiplier_10ccs_49_io_in_a),
    .io_in_b(FP_multiplier_10ccs_49_io_in_b),
    .io_out_s(FP_multiplier_10ccs_49_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_50 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_50_clock),
    .reset(FP_multiplier_10ccs_50_reset),
    .io_in_en(FP_multiplier_10ccs_50_io_in_en),
    .io_in_a(FP_multiplier_10ccs_50_io_in_a),
    .io_in_b(FP_multiplier_10ccs_50_io_in_b),
    .io_out_s(FP_multiplier_10ccs_50_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_51 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_51_clock),
    .reset(FP_multiplier_10ccs_51_reset),
    .io_in_en(FP_multiplier_10ccs_51_io_in_en),
    .io_in_a(FP_multiplier_10ccs_51_io_in_a),
    .io_in_b(FP_multiplier_10ccs_51_io_in_b),
    .io_out_s(FP_multiplier_10ccs_51_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_52 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_52_clock),
    .reset(FP_multiplier_10ccs_52_reset),
    .io_in_en(FP_multiplier_10ccs_52_io_in_en),
    .io_in_a(FP_multiplier_10ccs_52_io_in_a),
    .io_in_b(FP_multiplier_10ccs_52_io_in_b),
    .io_out_s(FP_multiplier_10ccs_52_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_53 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_53_clock),
    .reset(FP_multiplier_10ccs_53_reset),
    .io_in_en(FP_multiplier_10ccs_53_io_in_en),
    .io_in_a(FP_multiplier_10ccs_53_io_in_a),
    .io_in_b(FP_multiplier_10ccs_53_io_in_b),
    .io_out_s(FP_multiplier_10ccs_53_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_54 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_54_clock),
    .reset(FP_multiplier_10ccs_54_reset),
    .io_in_en(FP_multiplier_10ccs_54_io_in_en),
    .io_in_a(FP_multiplier_10ccs_54_io_in_a),
    .io_in_b(FP_multiplier_10ccs_54_io_in_b),
    .io_out_s(FP_multiplier_10ccs_54_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_55 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_55_clock),
    .reset(FP_multiplier_10ccs_55_reset),
    .io_in_en(FP_multiplier_10ccs_55_io_in_en),
    .io_in_a(FP_multiplier_10ccs_55_io_in_a),
    .io_in_b(FP_multiplier_10ccs_55_io_in_b),
    .io_out_s(FP_multiplier_10ccs_55_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_56 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_56_clock),
    .reset(FP_multiplier_10ccs_56_reset),
    .io_in_en(FP_multiplier_10ccs_56_io_in_en),
    .io_in_a(FP_multiplier_10ccs_56_io_in_a),
    .io_in_b(FP_multiplier_10ccs_56_io_in_b),
    .io_out_s(FP_multiplier_10ccs_56_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_57 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_57_clock),
    .reset(FP_multiplier_10ccs_57_reset),
    .io_in_en(FP_multiplier_10ccs_57_io_in_en),
    .io_in_a(FP_multiplier_10ccs_57_io_in_a),
    .io_in_b(FP_multiplier_10ccs_57_io_in_b),
    .io_out_s(FP_multiplier_10ccs_57_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_58 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_58_clock),
    .reset(FP_multiplier_10ccs_58_reset),
    .io_in_en(FP_multiplier_10ccs_58_io_in_en),
    .io_in_a(FP_multiplier_10ccs_58_io_in_a),
    .io_in_b(FP_multiplier_10ccs_58_io_in_b),
    .io_out_s(FP_multiplier_10ccs_58_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_59 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_59_clock),
    .reset(FP_multiplier_10ccs_59_reset),
    .io_in_en(FP_multiplier_10ccs_59_io_in_en),
    .io_in_a(FP_multiplier_10ccs_59_io_in_a),
    .io_in_b(FP_multiplier_10ccs_59_io_in_b),
    .io_out_s(FP_multiplier_10ccs_59_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_60 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_60_clock),
    .reset(FP_multiplier_10ccs_60_reset),
    .io_in_en(FP_multiplier_10ccs_60_io_in_en),
    .io_in_a(FP_multiplier_10ccs_60_io_in_a),
    .io_in_b(FP_multiplier_10ccs_60_io_in_b),
    .io_out_s(FP_multiplier_10ccs_60_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_61 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_61_clock),
    .reset(FP_multiplier_10ccs_61_reset),
    .io_in_en(FP_multiplier_10ccs_61_io_in_en),
    .io_in_a(FP_multiplier_10ccs_61_io_in_a),
    .io_in_b(FP_multiplier_10ccs_61_io_in_b),
    .io_out_s(FP_multiplier_10ccs_61_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_62 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_62_clock),
    .reset(FP_multiplier_10ccs_62_reset),
    .io_in_en(FP_multiplier_10ccs_62_io_in_en),
    .io_in_a(FP_multiplier_10ccs_62_io_in_a),
    .io_in_b(FP_multiplier_10ccs_62_io_in_b),
    .io_out_s(FP_multiplier_10ccs_62_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_63 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_63_clock),
    .reset(FP_multiplier_10ccs_63_reset),
    .io_in_en(FP_multiplier_10ccs_63_io_in_en),
    .io_in_a(FP_multiplier_10ccs_63_io_in_a),
    .io_in_b(FP_multiplier_10ccs_63_io_in_b),
    .io_out_s(FP_multiplier_10ccs_63_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_64 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_64_clock),
    .reset(FP_multiplier_10ccs_64_reset),
    .io_in_en(FP_multiplier_10ccs_64_io_in_en),
    .io_in_a(FP_multiplier_10ccs_64_io_in_a),
    .io_in_b(FP_multiplier_10ccs_64_io_in_b),
    .io_out_s(FP_multiplier_10ccs_64_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_65 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_65_clock),
    .reset(FP_multiplier_10ccs_65_reset),
    .io_in_en(FP_multiplier_10ccs_65_io_in_en),
    .io_in_a(FP_multiplier_10ccs_65_io_in_a),
    .io_in_b(FP_multiplier_10ccs_65_io_in_b),
    .io_out_s(FP_multiplier_10ccs_65_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_66 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_66_clock),
    .reset(FP_multiplier_10ccs_66_reset),
    .io_in_en(FP_multiplier_10ccs_66_io_in_en),
    .io_in_a(FP_multiplier_10ccs_66_io_in_a),
    .io_in_b(FP_multiplier_10ccs_66_io_in_b),
    .io_out_s(FP_multiplier_10ccs_66_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_67 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_67_clock),
    .reset(FP_multiplier_10ccs_67_reset),
    .io_in_en(FP_multiplier_10ccs_67_io_in_en),
    .io_in_a(FP_multiplier_10ccs_67_io_in_a),
    .io_in_b(FP_multiplier_10ccs_67_io_in_b),
    .io_out_s(FP_multiplier_10ccs_67_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_68 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_68_clock),
    .reset(FP_multiplier_10ccs_68_reset),
    .io_in_en(FP_multiplier_10ccs_68_io_in_en),
    .io_in_a(FP_multiplier_10ccs_68_io_in_a),
    .io_in_b(FP_multiplier_10ccs_68_io_in_b),
    .io_out_s(FP_multiplier_10ccs_68_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_69 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_69_clock),
    .reset(FP_multiplier_10ccs_69_reset),
    .io_in_en(FP_multiplier_10ccs_69_io_in_en),
    .io_in_a(FP_multiplier_10ccs_69_io_in_a),
    .io_in_b(FP_multiplier_10ccs_69_io_in_b),
    .io_out_s(FP_multiplier_10ccs_69_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_70 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_70_clock),
    .reset(FP_multiplier_10ccs_70_reset),
    .io_in_en(FP_multiplier_10ccs_70_io_in_en),
    .io_in_a(FP_multiplier_10ccs_70_io_in_a),
    .io_in_b(FP_multiplier_10ccs_70_io_in_b),
    .io_out_s(FP_multiplier_10ccs_70_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_71 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_71_clock),
    .reset(FP_multiplier_10ccs_71_reset),
    .io_in_en(FP_multiplier_10ccs_71_io_in_en),
    .io_in_a(FP_multiplier_10ccs_71_io_in_a),
    .io_in_b(FP_multiplier_10ccs_71_io_in_b),
    .io_out_s(FP_multiplier_10ccs_71_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_72 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_72_clock),
    .reset(FP_multiplier_10ccs_72_reset),
    .io_in_en(FP_multiplier_10ccs_72_io_in_en),
    .io_in_a(FP_multiplier_10ccs_72_io_in_a),
    .io_in_b(FP_multiplier_10ccs_72_io_in_b),
    .io_out_s(FP_multiplier_10ccs_72_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_73 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_73_clock),
    .reset(FP_multiplier_10ccs_73_reset),
    .io_in_en(FP_multiplier_10ccs_73_io_in_en),
    .io_in_a(FP_multiplier_10ccs_73_io_in_a),
    .io_in_b(FP_multiplier_10ccs_73_io_in_b),
    .io_out_s(FP_multiplier_10ccs_73_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_74 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_74_clock),
    .reset(FP_multiplier_10ccs_74_reset),
    .io_in_en(FP_multiplier_10ccs_74_io_in_en),
    .io_in_a(FP_multiplier_10ccs_74_io_in_a),
    .io_in_b(FP_multiplier_10ccs_74_io_in_b),
    .io_out_s(FP_multiplier_10ccs_74_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_75 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_75_clock),
    .reset(FP_multiplier_10ccs_75_reset),
    .io_in_en(FP_multiplier_10ccs_75_io_in_en),
    .io_in_a(FP_multiplier_10ccs_75_io_in_a),
    .io_in_b(FP_multiplier_10ccs_75_io_in_b),
    .io_out_s(FP_multiplier_10ccs_75_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_76 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_76_clock),
    .reset(FP_multiplier_10ccs_76_reset),
    .io_in_en(FP_multiplier_10ccs_76_io_in_en),
    .io_in_a(FP_multiplier_10ccs_76_io_in_a),
    .io_in_b(FP_multiplier_10ccs_76_io_in_b),
    .io_out_s(FP_multiplier_10ccs_76_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_77 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_77_clock),
    .reset(FP_multiplier_10ccs_77_reset),
    .io_in_en(FP_multiplier_10ccs_77_io_in_en),
    .io_in_a(FP_multiplier_10ccs_77_io_in_a),
    .io_in_b(FP_multiplier_10ccs_77_io_in_b),
    .io_out_s(FP_multiplier_10ccs_77_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_78 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_78_clock),
    .reset(FP_multiplier_10ccs_78_reset),
    .io_in_en(FP_multiplier_10ccs_78_io_in_en),
    .io_in_a(FP_multiplier_10ccs_78_io_in_a),
    .io_in_b(FP_multiplier_10ccs_78_io_in_b),
    .io_out_s(FP_multiplier_10ccs_78_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_79 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_79_clock),
    .reset(FP_multiplier_10ccs_79_reset),
    .io_in_en(FP_multiplier_10ccs_79_io_in_en),
    .io_in_a(FP_multiplier_10ccs_79_io_in_a),
    .io_in_b(FP_multiplier_10ccs_79_io_in_b),
    .io_out_s(FP_multiplier_10ccs_79_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_80 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_80_clock),
    .reset(FP_multiplier_10ccs_80_reset),
    .io_in_en(FP_multiplier_10ccs_80_io_in_en),
    .io_in_a(FP_multiplier_10ccs_80_io_in_a),
    .io_in_b(FP_multiplier_10ccs_80_io_in_b),
    .io_out_s(FP_multiplier_10ccs_80_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_81 ( // @[FloatingPointDesigns.scala 2206:69]
    .clock(FP_multiplier_10ccs_81_clock),
    .reset(FP_multiplier_10ccs_81_reset),
    .io_in_en(FP_multiplier_10ccs_81_io_in_en),
    .io_in_a(FP_multiplier_10ccs_81_io_in_a),
    .io_in_b(FP_multiplier_10ccs_81_io_in_b),
    .io_out_s(FP_multiplier_10ccs_81_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_16 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_16_clock),
    .reset(FP_subtractor_13ccs_16_reset),
    .io_in_en(FP_subtractor_13ccs_16_io_in_en),
    .io_in_a(FP_subtractor_13ccs_16_io_in_a),
    .io_in_b(FP_subtractor_13ccs_16_io_in_b),
    .io_out_s(FP_subtractor_13ccs_16_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_17 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_17_clock),
    .reset(FP_subtractor_13ccs_17_reset),
    .io_in_en(FP_subtractor_13ccs_17_io_in_en),
    .io_in_a(FP_subtractor_13ccs_17_io_in_a),
    .io_in_b(FP_subtractor_13ccs_17_io_in_b),
    .io_out_s(FP_subtractor_13ccs_17_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_18 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_18_clock),
    .reset(FP_subtractor_13ccs_18_reset),
    .io_in_en(FP_subtractor_13ccs_18_io_in_en),
    .io_in_a(FP_subtractor_13ccs_18_io_in_a),
    .io_in_b(FP_subtractor_13ccs_18_io_in_b),
    .io_out_s(FP_subtractor_13ccs_18_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_19 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_19_clock),
    .reset(FP_subtractor_13ccs_19_reset),
    .io_in_en(FP_subtractor_13ccs_19_io_in_en),
    .io_in_a(FP_subtractor_13ccs_19_io_in_a),
    .io_in_b(FP_subtractor_13ccs_19_io_in_b),
    .io_out_s(FP_subtractor_13ccs_19_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_20 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_20_clock),
    .reset(FP_subtractor_13ccs_20_reset),
    .io_in_en(FP_subtractor_13ccs_20_io_in_en),
    .io_in_a(FP_subtractor_13ccs_20_io_in_a),
    .io_in_b(FP_subtractor_13ccs_20_io_in_b),
    .io_out_s(FP_subtractor_13ccs_20_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_21 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_21_clock),
    .reset(FP_subtractor_13ccs_21_reset),
    .io_in_en(FP_subtractor_13ccs_21_io_in_en),
    .io_in_a(FP_subtractor_13ccs_21_io_in_a),
    .io_in_b(FP_subtractor_13ccs_21_io_in_b),
    .io_out_s(FP_subtractor_13ccs_21_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_22 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_22_clock),
    .reset(FP_subtractor_13ccs_22_reset),
    .io_in_en(FP_subtractor_13ccs_22_io_in_en),
    .io_in_a(FP_subtractor_13ccs_22_io_in_a),
    .io_in_b(FP_subtractor_13ccs_22_io_in_b),
    .io_out_s(FP_subtractor_13ccs_22_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_23 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_23_clock),
    .reset(FP_subtractor_13ccs_23_reset),
    .io_in_en(FP_subtractor_13ccs_23_io_in_en),
    .io_in_a(FP_subtractor_13ccs_23_io_in_a),
    .io_in_b(FP_subtractor_13ccs_23_io_in_b),
    .io_out_s(FP_subtractor_13ccs_23_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_24 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_24_clock),
    .reset(FP_subtractor_13ccs_24_reset),
    .io_in_en(FP_subtractor_13ccs_24_io_in_en),
    .io_in_a(FP_subtractor_13ccs_24_io_in_a),
    .io_in_b(FP_subtractor_13ccs_24_io_in_b),
    .io_out_s(FP_subtractor_13ccs_24_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_25 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_25_clock),
    .reset(FP_subtractor_13ccs_25_reset),
    .io_in_en(FP_subtractor_13ccs_25_io_in_en),
    .io_in_a(FP_subtractor_13ccs_25_io_in_a),
    .io_in_b(FP_subtractor_13ccs_25_io_in_b),
    .io_out_s(FP_subtractor_13ccs_25_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_26 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_26_clock),
    .reset(FP_subtractor_13ccs_26_reset),
    .io_in_en(FP_subtractor_13ccs_26_io_in_en),
    .io_in_a(FP_subtractor_13ccs_26_io_in_a),
    .io_in_b(FP_subtractor_13ccs_26_io_in_b),
    .io_out_s(FP_subtractor_13ccs_26_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_27 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_27_clock),
    .reset(FP_subtractor_13ccs_27_reset),
    .io_in_en(FP_subtractor_13ccs_27_io_in_en),
    .io_in_a(FP_subtractor_13ccs_27_io_in_a),
    .io_in_b(FP_subtractor_13ccs_27_io_in_b),
    .io_out_s(FP_subtractor_13ccs_27_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_28 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_28_clock),
    .reset(FP_subtractor_13ccs_28_reset),
    .io_in_en(FP_subtractor_13ccs_28_io_in_en),
    .io_in_a(FP_subtractor_13ccs_28_io_in_a),
    .io_in_b(FP_subtractor_13ccs_28_io_in_b),
    .io_out_s(FP_subtractor_13ccs_28_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_29 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_29_clock),
    .reset(FP_subtractor_13ccs_29_reset),
    .io_in_en(FP_subtractor_13ccs_29_io_in_en),
    .io_in_a(FP_subtractor_13ccs_29_io_in_a),
    .io_in_b(FP_subtractor_13ccs_29_io_in_b),
    .io_out_s(FP_subtractor_13ccs_29_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_30 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_30_clock),
    .reset(FP_subtractor_13ccs_30_reset),
    .io_in_en(FP_subtractor_13ccs_30_io_in_en),
    .io_in_a(FP_subtractor_13ccs_30_io_in_a),
    .io_in_b(FP_subtractor_13ccs_30_io_in_b),
    .io_out_s(FP_subtractor_13ccs_30_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_31 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_31_clock),
    .reset(FP_subtractor_13ccs_31_reset),
    .io_in_en(FP_subtractor_13ccs_31_io_in_en),
    .io_in_a(FP_subtractor_13ccs_31_io_in_a),
    .io_in_b(FP_subtractor_13ccs_31_io_in_b),
    .io_out_s(FP_subtractor_13ccs_31_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_32 ( // @[FloatingPointDesigns.scala 2207:54]
    .clock(FP_subtractor_13ccs_32_clock),
    .reset(FP_subtractor_13ccs_32_reset),
    .io_in_en(FP_subtractor_13ccs_32_io_in_en),
    .io_in_a(FP_subtractor_13ccs_32_io_in_a),
    .io_in_b(FP_subtractor_13ccs_32_io_in_b),
    .io_out_s(FP_subtractor_13ccs_32_io_out_s)
  );
  assign io_out_s = {stage3_regs_r_16_1_8[31],FP_multiplier_10ccs_81_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2263:58]
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_io_in_a = {1'h0,result[30:0]}; // @[FloatingPointDesigns.scala 2143:48]
  assign FP_multiplier_10ccs_io_in_b = {1'h0,result[30:0]}; // @[FloatingPointDesigns.scala 2144:48]
  assign FP_multiplier_10ccs_1_clock = clock;
  assign FP_multiplier_10ccs_1_reset = reset;
  assign FP_multiplier_10ccs_1_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_1_io_in_a = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_1_io_in_b = {1'h0,stage1_regs_0_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_2_clock = clock;
  assign FP_multiplier_10ccs_2_reset = reset;
  assign FP_multiplier_10ccs_2_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_2_io_in_a = {1'h0,stage3_regs_0_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_2_io_in_b = FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_3_clock = clock;
  assign FP_multiplier_10ccs_3_reset = reset;
  assign FP_multiplier_10ccs_3_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_3_io_in_a = {1'h0,FP_multiplier_10ccs_2_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_3_io_in_b = {1'h0,FP_multiplier_10ccs_2_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_4_clock = clock;
  assign FP_multiplier_10ccs_4_reset = reset;
  assign FP_multiplier_10ccs_4_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_4_io_in_a = FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_4_io_in_b = {1'h0,stage1_regs_1_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_5_clock = clock;
  assign FP_multiplier_10ccs_5_reset = reset;
  assign FP_multiplier_10ccs_5_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_5_io_in_a = {1'h0,stage3_regs_1_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_5_io_in_b = FP_subtractor_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_6_clock = clock;
  assign FP_multiplier_10ccs_6_reset = reset;
  assign FP_multiplier_10ccs_6_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_6_io_in_a = {1'h0,FP_multiplier_10ccs_5_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_6_io_in_b = {1'h0,FP_multiplier_10ccs_5_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_7_clock = clock;
  assign FP_multiplier_10ccs_7_reset = reset;
  assign FP_multiplier_10ccs_7_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_7_io_in_a = FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_7_io_in_b = {1'h0,stage1_regs_2_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_8_clock = clock;
  assign FP_multiplier_10ccs_8_reset = reset;
  assign FP_multiplier_10ccs_8_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_8_io_in_a = {1'h0,stage3_regs_2_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_8_io_in_b = FP_subtractor_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_9_clock = clock;
  assign FP_multiplier_10ccs_9_reset = reset;
  assign FP_multiplier_10ccs_9_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_9_io_in_a = {1'h0,FP_multiplier_10ccs_8_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_9_io_in_b = {1'h0,FP_multiplier_10ccs_8_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_10_clock = clock;
  assign FP_multiplier_10ccs_10_reset = reset;
  assign FP_multiplier_10ccs_10_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_10_io_in_a = FP_multiplier_10ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_10_io_in_b = {1'h0,stage1_regs_3_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_11_clock = clock;
  assign FP_multiplier_10ccs_11_reset = reset;
  assign FP_multiplier_10ccs_11_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_11_io_in_a = {1'h0,stage3_regs_3_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_11_io_in_b = FP_subtractor_13ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_12_clock = clock;
  assign FP_multiplier_10ccs_12_reset = reset;
  assign FP_multiplier_10ccs_12_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_12_io_in_a = {1'h0,FP_multiplier_10ccs_11_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_12_io_in_b = {1'h0,FP_multiplier_10ccs_11_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_13_clock = clock;
  assign FP_multiplier_10ccs_13_reset = reset;
  assign FP_multiplier_10ccs_13_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_13_io_in_a = FP_multiplier_10ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_13_io_in_b = {1'h0,stage1_regs_4_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_14_clock = clock;
  assign FP_multiplier_10ccs_14_reset = reset;
  assign FP_multiplier_10ccs_14_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_14_io_in_a = {1'h0,stage3_regs_4_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_14_io_in_b = FP_subtractor_13ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_15_clock = clock;
  assign FP_multiplier_10ccs_15_reset = reset;
  assign FP_multiplier_10ccs_15_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_15_io_in_a = {1'h0,FP_multiplier_10ccs_14_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_15_io_in_b = {1'h0,FP_multiplier_10ccs_14_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_16_clock = clock;
  assign FP_multiplier_10ccs_16_reset = reset;
  assign FP_multiplier_10ccs_16_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_16_io_in_a = FP_multiplier_10ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_16_io_in_b = {1'h0,stage1_regs_5_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_17_clock = clock;
  assign FP_multiplier_10ccs_17_reset = reset;
  assign FP_multiplier_10ccs_17_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_17_io_in_a = {1'h0,stage3_regs_5_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_17_io_in_b = FP_subtractor_13ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_18_clock = clock;
  assign FP_multiplier_10ccs_18_reset = reset;
  assign FP_multiplier_10ccs_18_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_18_io_in_a = {1'h0,FP_multiplier_10ccs_17_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_18_io_in_b = {1'h0,FP_multiplier_10ccs_17_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_19_clock = clock;
  assign FP_multiplier_10ccs_19_reset = reset;
  assign FP_multiplier_10ccs_19_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_19_io_in_a = FP_multiplier_10ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_19_io_in_b = {1'h0,stage1_regs_6_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_20_clock = clock;
  assign FP_multiplier_10ccs_20_reset = reset;
  assign FP_multiplier_10ccs_20_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_20_io_in_a = {1'h0,stage3_regs_6_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_20_io_in_b = FP_subtractor_13ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_21_clock = clock;
  assign FP_multiplier_10ccs_21_reset = reset;
  assign FP_multiplier_10ccs_21_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_21_io_in_a = {1'h0,FP_multiplier_10ccs_20_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_21_io_in_b = {1'h0,FP_multiplier_10ccs_20_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_22_clock = clock;
  assign FP_multiplier_10ccs_22_reset = reset;
  assign FP_multiplier_10ccs_22_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_22_io_in_a = FP_multiplier_10ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_22_io_in_b = {1'h0,stage1_regs_7_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_23_clock = clock;
  assign FP_multiplier_10ccs_23_reset = reset;
  assign FP_multiplier_10ccs_23_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_23_io_in_a = {1'h0,stage3_regs_7_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_23_io_in_b = FP_subtractor_13ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_24_clock = clock;
  assign FP_multiplier_10ccs_24_reset = reset;
  assign FP_multiplier_10ccs_24_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_24_io_in_a = {1'h0,FP_multiplier_10ccs_23_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_24_io_in_b = {1'h0,FP_multiplier_10ccs_23_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_25_clock = clock;
  assign FP_multiplier_10ccs_25_reset = reset;
  assign FP_multiplier_10ccs_25_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_25_io_in_a = FP_multiplier_10ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_25_io_in_b = {1'h0,stage1_regs_8_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_26_clock = clock;
  assign FP_multiplier_10ccs_26_reset = reset;
  assign FP_multiplier_10ccs_26_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_26_io_in_a = {1'h0,stage3_regs_8_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_26_io_in_b = FP_subtractor_13ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_27_clock = clock;
  assign FP_multiplier_10ccs_27_reset = reset;
  assign FP_multiplier_10ccs_27_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_27_io_in_a = {1'h0,FP_multiplier_10ccs_26_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_27_io_in_b = {1'h0,FP_multiplier_10ccs_26_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_28_clock = clock;
  assign FP_multiplier_10ccs_28_reset = reset;
  assign FP_multiplier_10ccs_28_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_28_io_in_a = FP_multiplier_10ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_28_io_in_b = {1'h0,stage1_regs_9_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_29_clock = clock;
  assign FP_multiplier_10ccs_29_reset = reset;
  assign FP_multiplier_10ccs_29_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_29_io_in_a = {1'h0,stage3_regs_9_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_29_io_in_b = FP_subtractor_13ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_30_clock = clock;
  assign FP_multiplier_10ccs_30_reset = reset;
  assign FP_multiplier_10ccs_30_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_30_io_in_a = {1'h0,FP_multiplier_10ccs_29_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_30_io_in_b = {1'h0,FP_multiplier_10ccs_29_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_31_clock = clock;
  assign FP_multiplier_10ccs_31_reset = reset;
  assign FP_multiplier_10ccs_31_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_31_io_in_a = FP_multiplier_10ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_31_io_in_b = {1'h0,stage1_regs_10_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_32_clock = clock;
  assign FP_multiplier_10ccs_32_reset = reset;
  assign FP_multiplier_10ccs_32_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_32_io_in_a = {1'h0,stage3_regs_10_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_32_io_in_b = FP_subtractor_13ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_33_clock = clock;
  assign FP_multiplier_10ccs_33_reset = reset;
  assign FP_multiplier_10ccs_33_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_33_io_in_a = {1'h0,FP_multiplier_10ccs_32_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_33_io_in_b = {1'h0,FP_multiplier_10ccs_32_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_34_clock = clock;
  assign FP_multiplier_10ccs_34_reset = reset;
  assign FP_multiplier_10ccs_34_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_34_io_in_a = FP_multiplier_10ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_34_io_in_b = {1'h0,stage1_regs_11_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_35_clock = clock;
  assign FP_multiplier_10ccs_35_reset = reset;
  assign FP_multiplier_10ccs_35_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_35_io_in_a = {1'h0,stage3_regs_11_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_35_io_in_b = FP_subtractor_13ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_36_clock = clock;
  assign FP_multiplier_10ccs_36_reset = reset;
  assign FP_multiplier_10ccs_36_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_36_io_in_a = {1'h0,FP_multiplier_10ccs_35_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_36_io_in_b = {1'h0,FP_multiplier_10ccs_35_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_37_clock = clock;
  assign FP_multiplier_10ccs_37_reset = reset;
  assign FP_multiplier_10ccs_37_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_37_io_in_a = FP_multiplier_10ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_37_io_in_b = {1'h0,stage1_regs_12_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_38_clock = clock;
  assign FP_multiplier_10ccs_38_reset = reset;
  assign FP_multiplier_10ccs_38_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_38_io_in_a = {1'h0,stage3_regs_12_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_38_io_in_b = FP_subtractor_13ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_39_clock = clock;
  assign FP_multiplier_10ccs_39_reset = reset;
  assign FP_multiplier_10ccs_39_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_39_io_in_a = {1'h0,FP_multiplier_10ccs_38_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_39_io_in_b = {1'h0,FP_multiplier_10ccs_38_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_40_clock = clock;
  assign FP_multiplier_10ccs_40_reset = reset;
  assign FP_multiplier_10ccs_40_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_40_io_in_a = FP_multiplier_10ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_40_io_in_b = {1'h0,stage1_regs_13_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_41_clock = clock;
  assign FP_multiplier_10ccs_41_reset = reset;
  assign FP_multiplier_10ccs_41_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_41_io_in_a = {1'h0,stage3_regs_13_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_41_io_in_b = FP_subtractor_13ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_42_clock = clock;
  assign FP_multiplier_10ccs_42_reset = reset;
  assign FP_multiplier_10ccs_42_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_42_io_in_a = {1'h0,FP_multiplier_10ccs_41_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_42_io_in_b = {1'h0,FP_multiplier_10ccs_41_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_43_clock = clock;
  assign FP_multiplier_10ccs_43_reset = reset;
  assign FP_multiplier_10ccs_43_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_43_io_in_a = FP_multiplier_10ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_43_io_in_b = {1'h0,stage1_regs_14_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_44_clock = clock;
  assign FP_multiplier_10ccs_44_reset = reset;
  assign FP_multiplier_10ccs_44_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_44_io_in_a = {1'h0,stage3_regs_14_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_44_io_in_b = FP_subtractor_13ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_multiplier_10ccs_45_clock = clock;
  assign FP_multiplier_10ccs_45_reset = reset;
  assign FP_multiplier_10ccs_45_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_45_io_in_a = {1'h0,FP_multiplier_10ccs_44_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2152:48]
  assign FP_multiplier_10ccs_45_io_in_b = {1'h0,FP_multiplier_10ccs_44_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2153:48]
  assign FP_multiplier_10ccs_46_clock = clock;
  assign FP_multiplier_10ccs_46_reset = reset;
  assign FP_multiplier_10ccs_46_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_46_io_in_a = FP_multiplier_10ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2156:34]
  assign FP_multiplier_10ccs_46_io_in_b = {1'h0,stage1_regs_15_1_8[30:0]}; // @[FloatingPointDesigns.scala 2157:46]
  assign FP_multiplier_10ccs_47_clock = clock;
  assign FP_multiplier_10ccs_47_reset = reset;
  assign FP_multiplier_10ccs_47_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2116:41]
  assign FP_multiplier_10ccs_47_io_in_a = {1'h0,stage3_regs_15_0_11[30:0]}; // @[FloatingPointDesigns.scala 2174:46]
  assign FP_multiplier_10ccs_47_io_in_b = FP_subtractor_13ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2175:34]
  assign FP_subtractor_13ccs_clock = clock;
  assign FP_subtractor_13ccs_reset = reset;
  assign FP_subtractor_13ccs_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_io_in_b = FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_1_clock = clock;
  assign FP_subtractor_13ccs_1_reset = reset;
  assign FP_subtractor_13ccs_1_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_1_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_1_io_in_b = FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_2_clock = clock;
  assign FP_subtractor_13ccs_2_reset = reset;
  assign FP_subtractor_13ccs_2_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_2_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_2_io_in_b = FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_3_clock = clock;
  assign FP_subtractor_13ccs_3_reset = reset;
  assign FP_subtractor_13ccs_3_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_3_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_3_io_in_b = FP_multiplier_10ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_4_clock = clock;
  assign FP_subtractor_13ccs_4_reset = reset;
  assign FP_subtractor_13ccs_4_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_4_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_4_io_in_b = FP_multiplier_10ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_5_clock = clock;
  assign FP_subtractor_13ccs_5_reset = reset;
  assign FP_subtractor_13ccs_5_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_5_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_5_io_in_b = FP_multiplier_10ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_6_clock = clock;
  assign FP_subtractor_13ccs_6_reset = reset;
  assign FP_subtractor_13ccs_6_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_6_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_6_io_in_b = FP_multiplier_10ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_7_clock = clock;
  assign FP_subtractor_13ccs_7_reset = reset;
  assign FP_subtractor_13ccs_7_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_7_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_7_io_in_b = FP_multiplier_10ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_8_clock = clock;
  assign FP_subtractor_13ccs_8_reset = reset;
  assign FP_subtractor_13ccs_8_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_8_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_8_io_in_b = FP_multiplier_10ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_9_clock = clock;
  assign FP_subtractor_13ccs_9_reset = reset;
  assign FP_subtractor_13ccs_9_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_9_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_9_io_in_b = FP_multiplier_10ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_10_clock = clock;
  assign FP_subtractor_13ccs_10_reset = reset;
  assign FP_subtractor_13ccs_10_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_10_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_10_io_in_b = FP_multiplier_10ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_11_clock = clock;
  assign FP_subtractor_13ccs_11_reset = reset;
  assign FP_subtractor_13ccs_11_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_11_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_11_io_in_b = FP_multiplier_10ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_12_clock = clock;
  assign FP_subtractor_13ccs_12_reset = reset;
  assign FP_subtractor_13ccs_12_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_12_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_12_io_in_b = FP_multiplier_10ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_13_clock = clock;
  assign FP_subtractor_13ccs_13_reset = reset;
  assign FP_subtractor_13ccs_13_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_13_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_13_io_in_b = FP_multiplier_10ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_14_clock = clock;
  assign FP_subtractor_13ccs_14_reset = reset;
  assign FP_subtractor_13ccs_14_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_14_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_14_io_in_b = FP_multiplier_10ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign FP_subtractor_13ccs_15_clock = clock;
  assign FP_subtractor_13ccs_15_reset = reset;
  assign FP_subtractor_13ccs_15_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2117:32]
  assign FP_subtractor_13ccs_15_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 2092:26 2093:16]
  assign FP_subtractor_13ccs_15_io_in_b = FP_multiplier_10ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2166:31]
  assign multiplier4_clock = clock;
  assign multiplier4_reset = reset;
  assign multiplier4_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2195:26]
  assign multiplier4_io_in_a = {1'h0,FP_multiplier_10ccs_47_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2196:37]
  assign multiplier4_io_in_b = {1'h0,FP_multiplier_10ccs_47_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2197:37]
  assign FP_multiplier_10ccs_48_clock = clock;
  assign FP_multiplier_10ccs_48_reset = reset;
  assign FP_multiplier_10ccs_48_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_48_io_in_a = {1'h0,multiplier4_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2232:50]
  assign FP_multiplier_10ccs_48_io_in_b = {1'h0,transition_regs_8[30:0]}; // @[FloatingPointDesigns.scala 2233:50]
  assign FP_multiplier_10ccs_49_clock = clock;
  assign FP_multiplier_10ccs_49_reset = reset;
  assign FP_multiplier_10ccs_49_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_49_io_in_a = {1'h0,stage2_regs_r_0_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_49_io_in_b = FP_subtractor_13ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_50_clock = clock;
  assign FP_multiplier_10ccs_50_reset = reset;
  assign FP_multiplier_10ccs_50_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_50_io_in_a = {1'h0,FP_multiplier_10ccs_49_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_50_io_in_b = {1'h0,stage3_regs_r_0_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_51_clock = clock;
  assign FP_multiplier_10ccs_51_reset = reset;
  assign FP_multiplier_10ccs_51_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_51_io_in_a = {1'h0,stage2_regs_r_1_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_51_io_in_b = FP_subtractor_13ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_52_clock = clock;
  assign FP_multiplier_10ccs_52_reset = reset;
  assign FP_multiplier_10ccs_52_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_52_io_in_a = {1'h0,FP_multiplier_10ccs_51_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_52_io_in_b = {1'h0,stage3_regs_r_1_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_53_clock = clock;
  assign FP_multiplier_10ccs_53_reset = reset;
  assign FP_multiplier_10ccs_53_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_53_io_in_a = {1'h0,stage2_regs_r_2_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_53_io_in_b = FP_subtractor_13ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_54_clock = clock;
  assign FP_multiplier_10ccs_54_reset = reset;
  assign FP_multiplier_10ccs_54_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_54_io_in_a = {1'h0,FP_multiplier_10ccs_53_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_54_io_in_b = {1'h0,stage3_regs_r_2_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_55_clock = clock;
  assign FP_multiplier_10ccs_55_reset = reset;
  assign FP_multiplier_10ccs_55_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_55_io_in_a = {1'h0,stage2_regs_r_3_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_55_io_in_b = FP_subtractor_13ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_56_clock = clock;
  assign FP_multiplier_10ccs_56_reset = reset;
  assign FP_multiplier_10ccs_56_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_56_io_in_a = {1'h0,FP_multiplier_10ccs_55_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_56_io_in_b = {1'h0,stage3_regs_r_3_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_57_clock = clock;
  assign FP_multiplier_10ccs_57_reset = reset;
  assign FP_multiplier_10ccs_57_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_57_io_in_a = {1'h0,stage2_regs_r_4_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_57_io_in_b = FP_subtractor_13ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_58_clock = clock;
  assign FP_multiplier_10ccs_58_reset = reset;
  assign FP_multiplier_10ccs_58_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_58_io_in_a = {1'h0,FP_multiplier_10ccs_57_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_58_io_in_b = {1'h0,stage3_regs_r_4_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_59_clock = clock;
  assign FP_multiplier_10ccs_59_reset = reset;
  assign FP_multiplier_10ccs_59_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_59_io_in_a = {1'h0,stage2_regs_r_5_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_59_io_in_b = FP_subtractor_13ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_60_clock = clock;
  assign FP_multiplier_10ccs_60_reset = reset;
  assign FP_multiplier_10ccs_60_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_60_io_in_a = {1'h0,FP_multiplier_10ccs_59_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_60_io_in_b = {1'h0,stage3_regs_r_5_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_61_clock = clock;
  assign FP_multiplier_10ccs_61_reset = reset;
  assign FP_multiplier_10ccs_61_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_61_io_in_a = {1'h0,stage2_regs_r_6_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_61_io_in_b = FP_subtractor_13ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_62_clock = clock;
  assign FP_multiplier_10ccs_62_reset = reset;
  assign FP_multiplier_10ccs_62_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_62_io_in_a = {1'h0,FP_multiplier_10ccs_61_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_62_io_in_b = {1'h0,stage3_regs_r_6_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_63_clock = clock;
  assign FP_multiplier_10ccs_63_reset = reset;
  assign FP_multiplier_10ccs_63_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_63_io_in_a = {1'h0,stage2_regs_r_7_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_63_io_in_b = FP_subtractor_13ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_64_clock = clock;
  assign FP_multiplier_10ccs_64_reset = reset;
  assign FP_multiplier_10ccs_64_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_64_io_in_a = {1'h0,FP_multiplier_10ccs_63_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_64_io_in_b = {1'h0,stage3_regs_r_7_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_65_clock = clock;
  assign FP_multiplier_10ccs_65_reset = reset;
  assign FP_multiplier_10ccs_65_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_65_io_in_a = {1'h0,stage2_regs_r_8_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_65_io_in_b = FP_subtractor_13ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_66_clock = clock;
  assign FP_multiplier_10ccs_66_reset = reset;
  assign FP_multiplier_10ccs_66_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_66_io_in_a = {1'h0,FP_multiplier_10ccs_65_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_66_io_in_b = {1'h0,stage3_regs_r_8_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_67_clock = clock;
  assign FP_multiplier_10ccs_67_reset = reset;
  assign FP_multiplier_10ccs_67_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_67_io_in_a = {1'h0,stage2_regs_r_9_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_67_io_in_b = FP_subtractor_13ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_68_clock = clock;
  assign FP_multiplier_10ccs_68_reset = reset;
  assign FP_multiplier_10ccs_68_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_68_io_in_a = {1'h0,FP_multiplier_10ccs_67_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_68_io_in_b = {1'h0,stage3_regs_r_9_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_69_clock = clock;
  assign FP_multiplier_10ccs_69_reset = reset;
  assign FP_multiplier_10ccs_69_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_69_io_in_a = {1'h0,stage2_regs_r_10_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_69_io_in_b = FP_subtractor_13ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_70_clock = clock;
  assign FP_multiplier_10ccs_70_reset = reset;
  assign FP_multiplier_10ccs_70_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_70_io_in_a = {1'h0,FP_multiplier_10ccs_69_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_70_io_in_b = {1'h0,stage3_regs_r_10_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_71_clock = clock;
  assign FP_multiplier_10ccs_71_reset = reset;
  assign FP_multiplier_10ccs_71_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_71_io_in_a = {1'h0,stage2_regs_r_11_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_71_io_in_b = FP_subtractor_13ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_72_clock = clock;
  assign FP_multiplier_10ccs_72_reset = reset;
  assign FP_multiplier_10ccs_72_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_72_io_in_a = {1'h0,FP_multiplier_10ccs_71_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_72_io_in_b = {1'h0,stage3_regs_r_11_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_73_clock = clock;
  assign FP_multiplier_10ccs_73_reset = reset;
  assign FP_multiplier_10ccs_73_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_73_io_in_a = {1'h0,stage2_regs_r_12_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_73_io_in_b = FP_subtractor_13ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_74_clock = clock;
  assign FP_multiplier_10ccs_74_reset = reset;
  assign FP_multiplier_10ccs_74_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_74_io_in_a = {1'h0,FP_multiplier_10ccs_73_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_74_io_in_b = {1'h0,stage3_regs_r_12_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_75_clock = clock;
  assign FP_multiplier_10ccs_75_reset = reset;
  assign FP_multiplier_10ccs_75_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_75_io_in_a = {1'h0,stage2_regs_r_13_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_75_io_in_b = FP_subtractor_13ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_76_clock = clock;
  assign FP_multiplier_10ccs_76_reset = reset;
  assign FP_multiplier_10ccs_76_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_76_io_in_a = {1'h0,FP_multiplier_10ccs_75_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_76_io_in_b = {1'h0,stage3_regs_r_13_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_77_clock = clock;
  assign FP_multiplier_10ccs_77_reset = reset;
  assign FP_multiplier_10ccs_77_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_77_io_in_a = {1'h0,stage2_regs_r_14_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_77_io_in_b = FP_subtractor_13ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_78_clock = clock;
  assign FP_multiplier_10ccs_78_reset = reset;
  assign FP_multiplier_10ccs_78_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_78_io_in_a = {1'h0,FP_multiplier_10ccs_77_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_78_io_in_b = {1'h0,stage3_regs_r_14_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_79_clock = clock;
  assign FP_multiplier_10ccs_79_reset = reset;
  assign FP_multiplier_10ccs_79_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_79_io_in_a = {1'h0,stage2_regs_r_15_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_79_io_in_b = FP_subtractor_13ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_multiplier_10ccs_80_clock = clock;
  assign FP_multiplier_10ccs_80_reset = reset;
  assign FP_multiplier_10ccs_80_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_80_io_in_a = {1'h0,FP_multiplier_10ccs_79_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2241:50]
  assign FP_multiplier_10ccs_80_io_in_b = {1'h0,stage3_regs_r_15_1_8[30:0]}; // @[FloatingPointDesigns.scala 2242:50]
  assign FP_multiplier_10ccs_81_clock = clock;
  assign FP_multiplier_10ccs_81_reset = reset;
  assign FP_multiplier_10ccs_81_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2208:43]
  assign FP_multiplier_10ccs_81_io_in_a = {1'h0,stage2_regs_r_16_0_11[30:0]}; // @[FloatingPointDesigns.scala 2254:48]
  assign FP_multiplier_10ccs_81_io_in_b = FP_subtractor_13ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2255:36]
  assign FP_subtractor_13ccs_16_clock = clock;
  assign FP_subtractor_13ccs_16_reset = reset;
  assign FP_subtractor_13ccs_16_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_16_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_16_io_in_b = FP_multiplier_10ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_17_clock = clock;
  assign FP_subtractor_13ccs_17_reset = reset;
  assign FP_subtractor_13ccs_17_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_17_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_17_io_in_b = FP_multiplier_10ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_18_clock = clock;
  assign FP_subtractor_13ccs_18_reset = reset;
  assign FP_subtractor_13ccs_18_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_18_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_18_io_in_b = FP_multiplier_10ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_19_clock = clock;
  assign FP_subtractor_13ccs_19_reset = reset;
  assign FP_subtractor_13ccs_19_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_19_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_19_io_in_b = FP_multiplier_10ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_20_clock = clock;
  assign FP_subtractor_13ccs_20_reset = reset;
  assign FP_subtractor_13ccs_20_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_20_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_20_io_in_b = FP_multiplier_10ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_21_clock = clock;
  assign FP_subtractor_13ccs_21_reset = reset;
  assign FP_subtractor_13ccs_21_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_21_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_21_io_in_b = FP_multiplier_10ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_22_clock = clock;
  assign FP_subtractor_13ccs_22_reset = reset;
  assign FP_subtractor_13ccs_22_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_22_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_22_io_in_b = FP_multiplier_10ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_23_clock = clock;
  assign FP_subtractor_13ccs_23_reset = reset;
  assign FP_subtractor_13ccs_23_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_23_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_23_io_in_b = FP_multiplier_10ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_24_clock = clock;
  assign FP_subtractor_13ccs_24_reset = reset;
  assign FP_subtractor_13ccs_24_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_24_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_24_io_in_b = FP_multiplier_10ccs_64_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_25_clock = clock;
  assign FP_subtractor_13ccs_25_reset = reset;
  assign FP_subtractor_13ccs_25_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_25_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_25_io_in_b = FP_multiplier_10ccs_66_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_26_clock = clock;
  assign FP_subtractor_13ccs_26_reset = reset;
  assign FP_subtractor_13ccs_26_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_26_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_26_io_in_b = FP_multiplier_10ccs_68_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_27_clock = clock;
  assign FP_subtractor_13ccs_27_reset = reset;
  assign FP_subtractor_13ccs_27_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_27_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_27_io_in_b = FP_multiplier_10ccs_70_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_28_clock = clock;
  assign FP_subtractor_13ccs_28_reset = reset;
  assign FP_subtractor_13ccs_28_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_28_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_28_io_in_b = FP_multiplier_10ccs_72_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_29_clock = clock;
  assign FP_subtractor_13ccs_29_reset = reset;
  assign FP_subtractor_13ccs_29_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_29_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_29_io_in_b = FP_multiplier_10ccs_74_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_30_clock = clock;
  assign FP_subtractor_13ccs_30_reset = reset;
  assign FP_subtractor_13ccs_30_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_30_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_30_io_in_b = FP_multiplier_10ccs_76_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_31_clock = clock;
  assign FP_subtractor_13ccs_31_reset = reset;
  assign FP_subtractor_13ccs_31_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_31_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_31_io_in_b = FP_multiplier_10ccs_78_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  assign FP_subtractor_13ccs_32_clock = clock;
  assign FP_subtractor_13ccs_32_reset = reset;
  assign FP_subtractor_13ccs_32_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2209:34]
  assign FP_subtractor_13ccs_32_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 2094:19 2095:9]
  assign FP_subtractor_13ccs_32_io_in_b = FP_multiplier_10ccs_80_io_out_s; // @[FloatingPointDesigns.scala 2246:33]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_0 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2137:28]
      x_n_0 <= result; // @[FloatingPointDesigns.scala 2138:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_1 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_1 <= stage1_regs_0_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_2 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_2 <= stage2_regs_0_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_4 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_4 <= FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_5 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_5 <= stage1_regs_1_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_6 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_6 <= stage2_regs_1_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_8 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_8 <= FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_9 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_9 <= stage1_regs_2_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_10 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_10 <= stage2_regs_2_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_12 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_12 <= FP_multiplier_10ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_13 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_13 <= stage1_regs_3_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_14 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_14 <= stage2_regs_3_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_16 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_16 <= FP_multiplier_10ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_17 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_17 <= stage1_regs_4_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_18 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_18 <= stage2_regs_4_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_20 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_20 <= FP_multiplier_10ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_21 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_21 <= stage1_regs_5_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_22 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_22 <= stage2_regs_5_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_24 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_24 <= FP_multiplier_10ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_25 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_25 <= stage1_regs_6_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_26 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_26 <= stage2_regs_6_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_28 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_28 <= FP_multiplier_10ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_29 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_29 <= stage1_regs_7_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_30 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_30 <= stage2_regs_7_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_32 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_32 <= FP_multiplier_10ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_33 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_33 <= stage1_regs_8_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_34 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_34 <= stage2_regs_8_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_36 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_36 <= FP_multiplier_10ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_37 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_37 <= stage1_regs_9_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_38 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_38 <= stage2_regs_9_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_40 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_40 <= FP_multiplier_10ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_41 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_41 <= stage1_regs_10_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_42 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_42 <= stage2_regs_10_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_44 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_44 <= FP_multiplier_10ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_45 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_45 <= stage1_regs_11_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_46 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_46 <= stage2_regs_11_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_48 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_48 <= FP_multiplier_10ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_49 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_49 <= stage1_regs_12_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_50 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_50 <= stage2_regs_12_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_52 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_52 <= FP_multiplier_10ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_53 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_53 <= stage1_regs_13_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_54 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_54 <= stage2_regs_13_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_56 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_56 <= FP_multiplier_10ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_57 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_57 <= stage1_regs_14_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_58 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_58 <= stage2_regs_14_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_60 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      x_n_60 <= FP_multiplier_10ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2147:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_61 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      x_n_61 <= stage1_regs_15_0_8; // @[FloatingPointDesigns.scala 2160:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2108:22]
      x_n_62 <= 32'h0; // @[FloatingPointDesigns.scala 2108:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      x_n_62 <= stage2_regs_15_0_8; // @[FloatingPointDesigns.scala 2169:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_0 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2137:28]
      a_2_0 <= _a_2_0_T_6; // @[FloatingPointDesigns.scala 2139:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_1 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_1 <= stage1_regs_0_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_2 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_2 <= stage2_regs_0_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_3 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_3 <= stage3_regs_0_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_4 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_4 <= stage4_regs_0_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_5 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_5 <= stage1_regs_1_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_6 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_6 <= stage2_regs_1_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_7 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_7 <= stage3_regs_1_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_8 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_8 <= stage4_regs_1_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_9 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_9 <= stage1_regs_2_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_10 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_10 <= stage2_regs_2_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_11 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_11 <= stage3_regs_2_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_12 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_12 <= stage4_regs_2_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_13 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_13 <= stage1_regs_3_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_14 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_14 <= stage2_regs_3_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_15 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_15 <= stage3_regs_3_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_16 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_16 <= stage4_regs_3_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_17 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_17 <= stage1_regs_4_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_18 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_18 <= stage2_regs_4_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_19 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_19 <= stage3_regs_4_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_20 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_20 <= stage4_regs_4_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_21 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_21 <= stage1_regs_5_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_22 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_22 <= stage2_regs_5_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_23 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_23 <= stage3_regs_5_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_24 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_24 <= stage4_regs_5_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_25 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_25 <= stage1_regs_6_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_26 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_26 <= stage2_regs_6_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_27 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_27 <= stage3_regs_6_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_28 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_28 <= stage4_regs_6_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_29 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_29 <= stage1_regs_7_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_30 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_30 <= stage2_regs_7_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_31 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_31 <= stage3_regs_7_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_32 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_32 <= stage4_regs_7_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_33 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_33 <= stage1_regs_8_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_34 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_34 <= stage2_regs_8_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_35 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_35 <= stage3_regs_8_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_36 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_36 <= stage4_regs_8_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_37 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_37 <= stage1_regs_9_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_38 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_38 <= stage2_regs_9_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_39 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_39 <= stage3_regs_9_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_40 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_40 <= stage4_regs_9_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_41 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_41 <= stage1_regs_10_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_42 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_42 <= stage2_regs_10_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_43 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_43 <= stage3_regs_10_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_44 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_44 <= stage4_regs_10_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_45 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_45 <= stage1_regs_11_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_46 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_46 <= stage2_regs_11_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_47 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_47 <= stage3_regs_11_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_48 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_48 <= stage4_regs_11_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_49 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_49 <= stage1_regs_12_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_50 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_50 <= stage2_regs_12_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_51 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_51 <= stage3_regs_12_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_52 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_52 <= stage4_regs_12_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_53 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_53 <= stage1_regs_13_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_54 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_54 <= stage2_regs_13_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_55 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_55 <= stage3_regs_13_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_56 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_56 <= stage4_regs_13_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_57 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_57 <= stage1_regs_14_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_58 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_58 <= stage2_regs_14_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_59 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_59 <= stage3_regs_14_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_60 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      a_2_60 <= stage4_regs_14_1_8; // @[FloatingPointDesigns.scala 2148:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_61 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      a_2_61 <= stage1_regs_15_1_8; // @[FloatingPointDesigns.scala 2159:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_62 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      a_2_62 <= stage2_regs_15_1_8; // @[FloatingPointDesigns.scala 2168:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2109:22]
      a_2_63 <= 32'h0; // @[FloatingPointDesigns.scala 2109:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      a_2_63 <= stage3_regs_15_1_11; // @[FloatingPointDesigns.scala 2177:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2137:28]
      stage1_regs_0_0_0 <= x_n_0; // @[FloatingPointDesigns.scala 2140:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_0_1 <= stage1_regs_0_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_0_2 <= stage1_regs_0_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_0_3 <= stage1_regs_0_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_0_4 <= stage1_regs_0_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_0_5 <= stage1_regs_0_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_0_6 <= stage1_regs_0_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_0_7 <= stage1_regs_0_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_0_8 <= stage1_regs_0_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2137:28]
      stage1_regs_0_1_0 <= a_2_0; // @[FloatingPointDesigns.scala 2141:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_1_1 <= stage1_regs_0_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_1_2 <= stage1_regs_0_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_1_3 <= stage1_regs_0_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_1_4 <= stage1_regs_0_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_1_5 <= stage1_regs_0_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_1_6 <= stage1_regs_0_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_1_7 <= stage1_regs_0_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_0_1_8 <= stage1_regs_0_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_1_0_0 <= x_n_4; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_0_1 <= stage1_regs_1_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_0_2 <= stage1_regs_1_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_0_3 <= stage1_regs_1_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_0_4 <= stage1_regs_1_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_0_5 <= stage1_regs_1_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_0_6 <= stage1_regs_1_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_0_7 <= stage1_regs_1_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_0_8 <= stage1_regs_1_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_1_1_0 <= a_2_4; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_1_1 <= stage1_regs_1_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_1_2 <= stage1_regs_1_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_1_3 <= stage1_regs_1_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_1_4 <= stage1_regs_1_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_1_5 <= stage1_regs_1_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_1_6 <= stage1_regs_1_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_1_7 <= stage1_regs_1_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_1_1_8 <= stage1_regs_1_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_2_0_0 <= x_n_8; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_0_1 <= stage1_regs_2_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_0_2 <= stage1_regs_2_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_0_3 <= stage1_regs_2_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_0_4 <= stage1_regs_2_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_0_5 <= stage1_regs_2_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_0_6 <= stage1_regs_2_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_0_7 <= stage1_regs_2_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_0_8 <= stage1_regs_2_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_2_1_0 <= a_2_8; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_1_1 <= stage1_regs_2_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_1_2 <= stage1_regs_2_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_1_3 <= stage1_regs_2_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_1_4 <= stage1_regs_2_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_1_5 <= stage1_regs_2_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_1_6 <= stage1_regs_2_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_1_7 <= stage1_regs_2_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_2_1_8 <= stage1_regs_2_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_3_0_0 <= x_n_12; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_0_1 <= stage1_regs_3_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_0_2 <= stage1_regs_3_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_0_3 <= stage1_regs_3_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_0_4 <= stage1_regs_3_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_0_5 <= stage1_regs_3_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_0_6 <= stage1_regs_3_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_0_7 <= stage1_regs_3_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_0_8 <= stage1_regs_3_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_3_1_0 <= a_2_12; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_1_1 <= stage1_regs_3_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_1_2 <= stage1_regs_3_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_1_3 <= stage1_regs_3_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_1_4 <= stage1_regs_3_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_1_5 <= stage1_regs_3_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_1_6 <= stage1_regs_3_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_1_7 <= stage1_regs_3_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_3_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_3_1_8 <= stage1_regs_3_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_4_0_0 <= x_n_16; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_0_1 <= stage1_regs_4_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_0_2 <= stage1_regs_4_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_0_3 <= stage1_regs_4_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_0_4 <= stage1_regs_4_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_0_5 <= stage1_regs_4_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_0_6 <= stage1_regs_4_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_0_7 <= stage1_regs_4_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_0_8 <= stage1_regs_4_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_4_1_0 <= a_2_16; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_1_1 <= stage1_regs_4_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_1_2 <= stage1_regs_4_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_1_3 <= stage1_regs_4_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_1_4 <= stage1_regs_4_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_1_5 <= stage1_regs_4_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_1_6 <= stage1_regs_4_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_1_7 <= stage1_regs_4_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_4_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_4_1_8 <= stage1_regs_4_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_5_0_0 <= x_n_20; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_0_1 <= stage1_regs_5_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_0_2 <= stage1_regs_5_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_0_3 <= stage1_regs_5_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_0_4 <= stage1_regs_5_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_0_5 <= stage1_regs_5_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_0_6 <= stage1_regs_5_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_0_7 <= stage1_regs_5_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_0_8 <= stage1_regs_5_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_5_1_0 <= a_2_20; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_1_1 <= stage1_regs_5_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_1_2 <= stage1_regs_5_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_1_3 <= stage1_regs_5_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_1_4 <= stage1_regs_5_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_1_5 <= stage1_regs_5_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_1_6 <= stage1_regs_5_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_1_7 <= stage1_regs_5_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_5_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_5_1_8 <= stage1_regs_5_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_6_0_0 <= x_n_24; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_0_1 <= stage1_regs_6_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_0_2 <= stage1_regs_6_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_0_3 <= stage1_regs_6_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_0_4 <= stage1_regs_6_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_0_5 <= stage1_regs_6_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_0_6 <= stage1_regs_6_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_0_7 <= stage1_regs_6_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_0_8 <= stage1_regs_6_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_6_1_0 <= a_2_24; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_1_1 <= stage1_regs_6_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_1_2 <= stage1_regs_6_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_1_3 <= stage1_regs_6_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_1_4 <= stage1_regs_6_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_1_5 <= stage1_regs_6_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_1_6 <= stage1_regs_6_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_1_7 <= stage1_regs_6_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_6_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_6_1_8 <= stage1_regs_6_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_7_0_0 <= x_n_28; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_0_1 <= stage1_regs_7_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_0_2 <= stage1_regs_7_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_0_3 <= stage1_regs_7_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_0_4 <= stage1_regs_7_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_0_5 <= stage1_regs_7_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_0_6 <= stage1_regs_7_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_0_7 <= stage1_regs_7_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_0_8 <= stage1_regs_7_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_7_1_0 <= a_2_28; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_1_1 <= stage1_regs_7_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_1_2 <= stage1_regs_7_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_1_3 <= stage1_regs_7_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_1_4 <= stage1_regs_7_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_1_5 <= stage1_regs_7_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_1_6 <= stage1_regs_7_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_1_7 <= stage1_regs_7_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_7_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_7_1_8 <= stage1_regs_7_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_8_0_0 <= x_n_32; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_0_1 <= stage1_regs_8_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_0_2 <= stage1_regs_8_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_0_3 <= stage1_regs_8_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_0_4 <= stage1_regs_8_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_0_5 <= stage1_regs_8_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_0_6 <= stage1_regs_8_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_0_7 <= stage1_regs_8_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_0_8 <= stage1_regs_8_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_8_1_0 <= a_2_32; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_1_1 <= stage1_regs_8_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_1_2 <= stage1_regs_8_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_1_3 <= stage1_regs_8_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_1_4 <= stage1_regs_8_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_1_5 <= stage1_regs_8_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_1_6 <= stage1_regs_8_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_1_7 <= stage1_regs_8_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_8_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_8_1_8 <= stage1_regs_8_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_9_0_0 <= x_n_36; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_0_1 <= stage1_regs_9_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_0_2 <= stage1_regs_9_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_0_3 <= stage1_regs_9_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_0_4 <= stage1_regs_9_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_0_5 <= stage1_regs_9_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_0_6 <= stage1_regs_9_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_0_7 <= stage1_regs_9_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_0_8 <= stage1_regs_9_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_9_1_0 <= a_2_36; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_1_1 <= stage1_regs_9_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_1_2 <= stage1_regs_9_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_1_3 <= stage1_regs_9_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_1_4 <= stage1_regs_9_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_1_5 <= stage1_regs_9_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_1_6 <= stage1_regs_9_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_1_7 <= stage1_regs_9_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_9_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_9_1_8 <= stage1_regs_9_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_10_0_0 <= x_n_40; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_0_1 <= stage1_regs_10_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_0_2 <= stage1_regs_10_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_0_3 <= stage1_regs_10_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_0_4 <= stage1_regs_10_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_0_5 <= stage1_regs_10_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_0_6 <= stage1_regs_10_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_0_7 <= stage1_regs_10_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_0_8 <= stage1_regs_10_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_10_1_0 <= a_2_40; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_1_1 <= stage1_regs_10_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_1_2 <= stage1_regs_10_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_1_3 <= stage1_regs_10_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_1_4 <= stage1_regs_10_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_1_5 <= stage1_regs_10_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_1_6 <= stage1_regs_10_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_1_7 <= stage1_regs_10_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_10_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_10_1_8 <= stage1_regs_10_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_11_0_0 <= x_n_44; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_0_1 <= stage1_regs_11_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_0_2 <= stage1_regs_11_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_0_3 <= stage1_regs_11_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_0_4 <= stage1_regs_11_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_0_5 <= stage1_regs_11_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_0_6 <= stage1_regs_11_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_0_7 <= stage1_regs_11_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_0_8 <= stage1_regs_11_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_11_1_0 <= a_2_44; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_1_1 <= stage1_regs_11_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_1_2 <= stage1_regs_11_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_1_3 <= stage1_regs_11_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_1_4 <= stage1_regs_11_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_1_5 <= stage1_regs_11_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_1_6 <= stage1_regs_11_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_1_7 <= stage1_regs_11_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_11_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_11_1_8 <= stage1_regs_11_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_12_0_0 <= x_n_48; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_0_1 <= stage1_regs_12_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_0_2 <= stage1_regs_12_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_0_3 <= stage1_regs_12_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_0_4 <= stage1_regs_12_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_0_5 <= stage1_regs_12_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_0_6 <= stage1_regs_12_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_0_7 <= stage1_regs_12_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_0_8 <= stage1_regs_12_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_12_1_0 <= a_2_48; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_1_1 <= stage1_regs_12_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_1_2 <= stage1_regs_12_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_1_3 <= stage1_regs_12_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_1_4 <= stage1_regs_12_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_1_5 <= stage1_regs_12_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_1_6 <= stage1_regs_12_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_1_7 <= stage1_regs_12_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_12_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_12_1_8 <= stage1_regs_12_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_13_0_0 <= x_n_52; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_0_1 <= stage1_regs_13_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_0_2 <= stage1_regs_13_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_0_3 <= stage1_regs_13_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_0_4 <= stage1_regs_13_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_0_5 <= stage1_regs_13_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_0_6 <= stage1_regs_13_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_0_7 <= stage1_regs_13_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_0_8 <= stage1_regs_13_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_13_1_0 <= a_2_52; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_1_1 <= stage1_regs_13_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_1_2 <= stage1_regs_13_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_1_3 <= stage1_regs_13_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_1_4 <= stage1_regs_13_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_1_5 <= stage1_regs_13_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_1_6 <= stage1_regs_13_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_1_7 <= stage1_regs_13_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_13_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_13_1_8 <= stage1_regs_13_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_14_0_0 <= x_n_56; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_0_1 <= stage1_regs_14_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_0_2 <= stage1_regs_14_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_0_3 <= stage1_regs_14_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_0_4 <= stage1_regs_14_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_0_5 <= stage1_regs_14_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_0_6 <= stage1_regs_14_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_0_7 <= stage1_regs_14_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_0_8 <= stage1_regs_14_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_14_1_0 <= a_2_56; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_1_1 <= stage1_regs_14_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_1_2 <= stage1_regs_14_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_1_3 <= stage1_regs_14_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_1_4 <= stage1_regs_14_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_1_5 <= stage1_regs_14_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_1_6 <= stage1_regs_14_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_1_7 <= stage1_regs_14_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_14_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_14_1_8 <= stage1_regs_14_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_15_0_0 <= x_n_60; // @[FloatingPointDesigns.scala 2149:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_0_1 <= stage1_regs_15_0_0; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_0_2 <= stage1_regs_15_0_1; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_0_3 <= stage1_regs_15_0_2; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_0_4 <= stage1_regs_15_0_3; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_0_5 <= stage1_regs_15_0_4; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_0_6 <= stage1_regs_15_0_5; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_0_7 <= stage1_regs_15_0_6; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_0_8 <= stage1_regs_15_0_7; // @[FloatingPointDesigns.scala 2126:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2146:28]
      stage1_regs_15_1_0 <= a_2_60; // @[FloatingPointDesigns.scala 2150:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_1_1 <= stage1_regs_15_1_0; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_1_2 <= stage1_regs_15_1_1; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_1_3 <= stage1_regs_15_1_2; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_1_4 <= stage1_regs_15_1_3; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_1_5 <= stage1_regs_15_1_4; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_1_6 <= stage1_regs_15_1_5; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_1_7 <= stage1_regs_15_1_6; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2110:30]
      stage1_regs_15_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2110:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage1_regs_15_1_8 <= stage1_regs_15_1_7; // @[FloatingPointDesigns.scala 2127:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_0_0_0 <= x_n_1; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_0_1 <= stage2_regs_0_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_0_2 <= stage2_regs_0_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_0_3 <= stage2_regs_0_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_0_4 <= stage2_regs_0_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_0_5 <= stage2_regs_0_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_0_6 <= stage2_regs_0_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_0_7 <= stage2_regs_0_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_0_8 <= stage2_regs_0_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_0_1_0 <= a_2_1; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_1_1 <= stage2_regs_0_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_1_2 <= stage2_regs_0_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_1_3 <= stage2_regs_0_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_1_4 <= stage2_regs_0_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_1_5 <= stage2_regs_0_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_1_6 <= stage2_regs_0_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_1_7 <= stage2_regs_0_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_0_1_8 <= stage2_regs_0_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_1_0_0 <= x_n_5; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_0_1 <= stage2_regs_1_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_0_2 <= stage2_regs_1_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_0_3 <= stage2_regs_1_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_0_4 <= stage2_regs_1_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_0_5 <= stage2_regs_1_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_0_6 <= stage2_regs_1_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_0_7 <= stage2_regs_1_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_0_8 <= stage2_regs_1_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_1_1_0 <= a_2_5; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_1_1 <= stage2_regs_1_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_1_2 <= stage2_regs_1_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_1_3 <= stage2_regs_1_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_1_4 <= stage2_regs_1_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_1_5 <= stage2_regs_1_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_1_6 <= stage2_regs_1_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_1_7 <= stage2_regs_1_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_1_1_8 <= stage2_regs_1_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_2_0_0 <= x_n_9; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_0_1 <= stage2_regs_2_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_0_2 <= stage2_regs_2_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_0_3 <= stage2_regs_2_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_0_4 <= stage2_regs_2_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_0_5 <= stage2_regs_2_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_0_6 <= stage2_regs_2_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_0_7 <= stage2_regs_2_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_0_8 <= stage2_regs_2_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_2_1_0 <= a_2_9; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_1_1 <= stage2_regs_2_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_1_2 <= stage2_regs_2_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_1_3 <= stage2_regs_2_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_1_4 <= stage2_regs_2_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_1_5 <= stage2_regs_2_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_1_6 <= stage2_regs_2_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_1_7 <= stage2_regs_2_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_2_1_8 <= stage2_regs_2_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_3_0_0 <= x_n_13; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_0_1 <= stage2_regs_3_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_0_2 <= stage2_regs_3_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_0_3 <= stage2_regs_3_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_0_4 <= stage2_regs_3_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_0_5 <= stage2_regs_3_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_0_6 <= stage2_regs_3_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_0_7 <= stage2_regs_3_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_0_8 <= stage2_regs_3_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_3_1_0 <= a_2_13; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_1_1 <= stage2_regs_3_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_1_2 <= stage2_regs_3_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_1_3 <= stage2_regs_3_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_1_4 <= stage2_regs_3_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_1_5 <= stage2_regs_3_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_1_6 <= stage2_regs_3_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_1_7 <= stage2_regs_3_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_3_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_3_1_8 <= stage2_regs_3_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_4_0_0 <= x_n_17; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_0_1 <= stage2_regs_4_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_0_2 <= stage2_regs_4_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_0_3 <= stage2_regs_4_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_0_4 <= stage2_regs_4_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_0_5 <= stage2_regs_4_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_0_6 <= stage2_regs_4_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_0_7 <= stage2_regs_4_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_0_8 <= stage2_regs_4_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_4_1_0 <= a_2_17; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_1_1 <= stage2_regs_4_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_1_2 <= stage2_regs_4_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_1_3 <= stage2_regs_4_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_1_4 <= stage2_regs_4_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_1_5 <= stage2_regs_4_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_1_6 <= stage2_regs_4_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_1_7 <= stage2_regs_4_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_4_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_4_1_8 <= stage2_regs_4_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_5_0_0 <= x_n_21; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_0_1 <= stage2_regs_5_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_0_2 <= stage2_regs_5_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_0_3 <= stage2_regs_5_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_0_4 <= stage2_regs_5_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_0_5 <= stage2_regs_5_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_0_6 <= stage2_regs_5_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_0_7 <= stage2_regs_5_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_0_8 <= stage2_regs_5_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_5_1_0 <= a_2_21; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_1_1 <= stage2_regs_5_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_1_2 <= stage2_regs_5_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_1_3 <= stage2_regs_5_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_1_4 <= stage2_regs_5_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_1_5 <= stage2_regs_5_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_1_6 <= stage2_regs_5_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_1_7 <= stage2_regs_5_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_5_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_5_1_8 <= stage2_regs_5_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_6_0_0 <= x_n_25; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_0_1 <= stage2_regs_6_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_0_2 <= stage2_regs_6_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_0_3 <= stage2_regs_6_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_0_4 <= stage2_regs_6_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_0_5 <= stage2_regs_6_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_0_6 <= stage2_regs_6_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_0_7 <= stage2_regs_6_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_0_8 <= stage2_regs_6_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_6_1_0 <= a_2_25; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_1_1 <= stage2_regs_6_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_1_2 <= stage2_regs_6_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_1_3 <= stage2_regs_6_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_1_4 <= stage2_regs_6_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_1_5 <= stage2_regs_6_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_1_6 <= stage2_regs_6_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_1_7 <= stage2_regs_6_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_6_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_6_1_8 <= stage2_regs_6_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_7_0_0 <= x_n_29; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_0_1 <= stage2_regs_7_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_0_2 <= stage2_regs_7_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_0_3 <= stage2_regs_7_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_0_4 <= stage2_regs_7_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_0_5 <= stage2_regs_7_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_0_6 <= stage2_regs_7_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_0_7 <= stage2_regs_7_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_0_8 <= stage2_regs_7_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_7_1_0 <= a_2_29; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_1_1 <= stage2_regs_7_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_1_2 <= stage2_regs_7_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_1_3 <= stage2_regs_7_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_1_4 <= stage2_regs_7_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_1_5 <= stage2_regs_7_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_1_6 <= stage2_regs_7_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_1_7 <= stage2_regs_7_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_7_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_7_1_8 <= stage2_regs_7_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_8_0_0 <= x_n_33; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_0_1 <= stage2_regs_8_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_0_2 <= stage2_regs_8_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_0_3 <= stage2_regs_8_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_0_4 <= stage2_regs_8_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_0_5 <= stage2_regs_8_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_0_6 <= stage2_regs_8_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_0_7 <= stage2_regs_8_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_0_8 <= stage2_regs_8_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_8_1_0 <= a_2_33; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_1_1 <= stage2_regs_8_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_1_2 <= stage2_regs_8_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_1_3 <= stage2_regs_8_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_1_4 <= stage2_regs_8_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_1_5 <= stage2_regs_8_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_1_6 <= stage2_regs_8_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_1_7 <= stage2_regs_8_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_8_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_8_1_8 <= stage2_regs_8_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_9_0_0 <= x_n_37; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_0_1 <= stage2_regs_9_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_0_2 <= stage2_regs_9_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_0_3 <= stage2_regs_9_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_0_4 <= stage2_regs_9_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_0_5 <= stage2_regs_9_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_0_6 <= stage2_regs_9_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_0_7 <= stage2_regs_9_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_0_8 <= stage2_regs_9_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_9_1_0 <= a_2_37; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_1_1 <= stage2_regs_9_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_1_2 <= stage2_regs_9_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_1_3 <= stage2_regs_9_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_1_4 <= stage2_regs_9_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_1_5 <= stage2_regs_9_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_1_6 <= stage2_regs_9_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_1_7 <= stage2_regs_9_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_9_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_9_1_8 <= stage2_regs_9_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_10_0_0 <= x_n_41; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_0_1 <= stage2_regs_10_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_0_2 <= stage2_regs_10_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_0_3 <= stage2_regs_10_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_0_4 <= stage2_regs_10_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_0_5 <= stage2_regs_10_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_0_6 <= stage2_regs_10_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_0_7 <= stage2_regs_10_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_0_8 <= stage2_regs_10_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_10_1_0 <= a_2_41; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_1_1 <= stage2_regs_10_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_1_2 <= stage2_regs_10_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_1_3 <= stage2_regs_10_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_1_4 <= stage2_regs_10_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_1_5 <= stage2_regs_10_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_1_6 <= stage2_regs_10_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_1_7 <= stage2_regs_10_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_10_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_10_1_8 <= stage2_regs_10_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_11_0_0 <= x_n_45; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_0_1 <= stage2_regs_11_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_0_2 <= stage2_regs_11_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_0_3 <= stage2_regs_11_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_0_4 <= stage2_regs_11_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_0_5 <= stage2_regs_11_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_0_6 <= stage2_regs_11_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_0_7 <= stage2_regs_11_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_0_8 <= stage2_regs_11_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_11_1_0 <= a_2_45; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_1_1 <= stage2_regs_11_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_1_2 <= stage2_regs_11_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_1_3 <= stage2_regs_11_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_1_4 <= stage2_regs_11_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_1_5 <= stage2_regs_11_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_1_6 <= stage2_regs_11_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_1_7 <= stage2_regs_11_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_11_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_11_1_8 <= stage2_regs_11_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_12_0_0 <= x_n_49; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_0_1 <= stage2_regs_12_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_0_2 <= stage2_regs_12_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_0_3 <= stage2_regs_12_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_0_4 <= stage2_regs_12_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_0_5 <= stage2_regs_12_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_0_6 <= stage2_regs_12_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_0_7 <= stage2_regs_12_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_0_8 <= stage2_regs_12_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_12_1_0 <= a_2_49; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_1_1 <= stage2_regs_12_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_1_2 <= stage2_regs_12_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_1_3 <= stage2_regs_12_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_1_4 <= stage2_regs_12_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_1_5 <= stage2_regs_12_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_1_6 <= stage2_regs_12_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_1_7 <= stage2_regs_12_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_12_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_12_1_8 <= stage2_regs_12_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_13_0_0 <= x_n_53; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_0_1 <= stage2_regs_13_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_0_2 <= stage2_regs_13_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_0_3 <= stage2_regs_13_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_0_4 <= stage2_regs_13_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_0_5 <= stage2_regs_13_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_0_6 <= stage2_regs_13_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_0_7 <= stage2_regs_13_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_0_8 <= stage2_regs_13_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_13_1_0 <= a_2_53; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_1_1 <= stage2_regs_13_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_1_2 <= stage2_regs_13_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_1_3 <= stage2_regs_13_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_1_4 <= stage2_regs_13_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_1_5 <= stage2_regs_13_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_1_6 <= stage2_regs_13_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_1_7 <= stage2_regs_13_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_13_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_13_1_8 <= stage2_regs_13_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_14_0_0 <= x_n_57; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_0_1 <= stage2_regs_14_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_0_2 <= stage2_regs_14_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_0_3 <= stage2_regs_14_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_0_4 <= stage2_regs_14_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_0_5 <= stage2_regs_14_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_0_6 <= stage2_regs_14_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_0_7 <= stage2_regs_14_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_0_8 <= stage2_regs_14_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_14_1_0 <= a_2_57; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_1_1 <= stage2_regs_14_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_1_2 <= stage2_regs_14_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_1_3 <= stage2_regs_14_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_1_4 <= stage2_regs_14_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_1_5 <= stage2_regs_14_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_1_6 <= stage2_regs_14_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_1_7 <= stage2_regs_14_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_14_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_14_1_8 <= stage2_regs_14_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_15_0_0 <= x_n_61; // @[FloatingPointDesigns.scala 2161:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_0_1 <= stage2_regs_15_0_0; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_0_2 <= stage2_regs_15_0_1; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_0_3 <= stage2_regs_15_0_2; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_0_4 <= stage2_regs_15_0_3; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_0_5 <= stage2_regs_15_0_4; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_0_6 <= stage2_regs_15_0_5; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_0_7 <= stage2_regs_15_0_6; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_0_8 <= stage2_regs_15_0_7; // @[FloatingPointDesigns.scala 2128:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2158:26]
      stage2_regs_15_1_0 <= a_2_61; // @[FloatingPointDesigns.scala 2162:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_1_1 <= stage2_regs_15_1_0; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_1_2 <= stage2_regs_15_1_1; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_1_3 <= stage2_regs_15_1_2; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_1_4 <= stage2_regs_15_1_3; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_1_5 <= stage2_regs_15_1_4; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_1_6 <= stage2_regs_15_1_5; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_1_7 <= stage2_regs_15_1_6; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2111:30]
      stage2_regs_15_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2111:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage2_regs_15_1_8 <= stage2_regs_15_1_7; // @[FloatingPointDesigns.scala 2129:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_0_0_0 <= x_n_2; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_0_1 <= stage3_regs_0_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_0_2 <= stage3_regs_0_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_0_3 <= stage3_regs_0_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_0_4 <= stage3_regs_0_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_0_5 <= stage3_regs_0_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_0_6 <= stage3_regs_0_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_0_7 <= stage3_regs_0_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_0_8 <= stage3_regs_0_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_0_9 <= stage3_regs_0_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_0_10 <= stage3_regs_0_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_0_11 <= stage3_regs_0_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_0_1_0 <= a_2_2; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_1_1 <= stage3_regs_0_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_1_2 <= stage3_regs_0_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_1_3 <= stage3_regs_0_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_1_4 <= stage3_regs_0_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_1_5 <= stage3_regs_0_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_1_6 <= stage3_regs_0_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_1_7 <= stage3_regs_0_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_1_8 <= stage3_regs_0_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_1_9 <= stage3_regs_0_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_1_10 <= stage3_regs_0_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_0_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_0_1_11 <= stage3_regs_0_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_1_0_0 <= x_n_6; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_0_1 <= stage3_regs_1_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_0_2 <= stage3_regs_1_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_0_3 <= stage3_regs_1_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_0_4 <= stage3_regs_1_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_0_5 <= stage3_regs_1_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_0_6 <= stage3_regs_1_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_0_7 <= stage3_regs_1_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_0_8 <= stage3_regs_1_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_0_9 <= stage3_regs_1_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_0_10 <= stage3_regs_1_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_0_11 <= stage3_regs_1_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_1_1_0 <= a_2_6; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_1_1 <= stage3_regs_1_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_1_2 <= stage3_regs_1_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_1_3 <= stage3_regs_1_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_1_4 <= stage3_regs_1_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_1_5 <= stage3_regs_1_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_1_6 <= stage3_regs_1_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_1_7 <= stage3_regs_1_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_1_8 <= stage3_regs_1_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_1_9 <= stage3_regs_1_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_1_10 <= stage3_regs_1_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_1_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_1_1_11 <= stage3_regs_1_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_2_0_0 <= x_n_10; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_0_1 <= stage3_regs_2_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_0_2 <= stage3_regs_2_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_0_3 <= stage3_regs_2_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_0_4 <= stage3_regs_2_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_0_5 <= stage3_regs_2_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_0_6 <= stage3_regs_2_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_0_7 <= stage3_regs_2_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_0_8 <= stage3_regs_2_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_0_9 <= stage3_regs_2_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_0_10 <= stage3_regs_2_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_0_11 <= stage3_regs_2_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_2_1_0 <= a_2_10; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_1_1 <= stage3_regs_2_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_1_2 <= stage3_regs_2_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_1_3 <= stage3_regs_2_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_1_4 <= stage3_regs_2_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_1_5 <= stage3_regs_2_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_1_6 <= stage3_regs_2_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_1_7 <= stage3_regs_2_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_1_8 <= stage3_regs_2_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_1_9 <= stage3_regs_2_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_1_10 <= stage3_regs_2_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_2_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_2_1_11 <= stage3_regs_2_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_3_0_0 <= x_n_14; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_0_1 <= stage3_regs_3_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_0_2 <= stage3_regs_3_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_0_3 <= stage3_regs_3_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_0_4 <= stage3_regs_3_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_0_5 <= stage3_regs_3_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_0_6 <= stage3_regs_3_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_0_7 <= stage3_regs_3_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_0_8 <= stage3_regs_3_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_0_9 <= stage3_regs_3_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_0_10 <= stage3_regs_3_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_0_11 <= stage3_regs_3_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_3_1_0 <= a_2_14; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_1_1 <= stage3_regs_3_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_1_2 <= stage3_regs_3_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_1_3 <= stage3_regs_3_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_1_4 <= stage3_regs_3_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_1_5 <= stage3_regs_3_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_1_6 <= stage3_regs_3_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_1_7 <= stage3_regs_3_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_1_8 <= stage3_regs_3_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_1_9 <= stage3_regs_3_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_1_10 <= stage3_regs_3_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_3_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_3_1_11 <= stage3_regs_3_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_4_0_0 <= x_n_18; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_0_1 <= stage3_regs_4_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_0_2 <= stage3_regs_4_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_0_3 <= stage3_regs_4_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_0_4 <= stage3_regs_4_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_0_5 <= stage3_regs_4_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_0_6 <= stage3_regs_4_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_0_7 <= stage3_regs_4_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_0_8 <= stage3_regs_4_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_0_9 <= stage3_regs_4_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_0_10 <= stage3_regs_4_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_0_11 <= stage3_regs_4_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_4_1_0 <= a_2_18; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_1_1 <= stage3_regs_4_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_1_2 <= stage3_regs_4_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_1_3 <= stage3_regs_4_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_1_4 <= stage3_regs_4_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_1_5 <= stage3_regs_4_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_1_6 <= stage3_regs_4_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_1_7 <= stage3_regs_4_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_1_8 <= stage3_regs_4_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_1_9 <= stage3_regs_4_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_1_10 <= stage3_regs_4_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_4_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_4_1_11 <= stage3_regs_4_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_5_0_0 <= x_n_22; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_0_1 <= stage3_regs_5_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_0_2 <= stage3_regs_5_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_0_3 <= stage3_regs_5_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_0_4 <= stage3_regs_5_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_0_5 <= stage3_regs_5_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_0_6 <= stage3_regs_5_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_0_7 <= stage3_regs_5_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_0_8 <= stage3_regs_5_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_0_9 <= stage3_regs_5_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_0_10 <= stage3_regs_5_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_0_11 <= stage3_regs_5_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_5_1_0 <= a_2_22; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_1_1 <= stage3_regs_5_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_1_2 <= stage3_regs_5_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_1_3 <= stage3_regs_5_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_1_4 <= stage3_regs_5_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_1_5 <= stage3_regs_5_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_1_6 <= stage3_regs_5_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_1_7 <= stage3_regs_5_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_1_8 <= stage3_regs_5_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_1_9 <= stage3_regs_5_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_1_10 <= stage3_regs_5_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_5_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_5_1_11 <= stage3_regs_5_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_6_0_0 <= x_n_26; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_0_1 <= stage3_regs_6_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_0_2 <= stage3_regs_6_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_0_3 <= stage3_regs_6_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_0_4 <= stage3_regs_6_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_0_5 <= stage3_regs_6_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_0_6 <= stage3_regs_6_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_0_7 <= stage3_regs_6_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_0_8 <= stage3_regs_6_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_0_9 <= stage3_regs_6_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_0_10 <= stage3_regs_6_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_0_11 <= stage3_regs_6_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_6_1_0 <= a_2_26; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_1_1 <= stage3_regs_6_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_1_2 <= stage3_regs_6_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_1_3 <= stage3_regs_6_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_1_4 <= stage3_regs_6_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_1_5 <= stage3_regs_6_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_1_6 <= stage3_regs_6_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_1_7 <= stage3_regs_6_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_1_8 <= stage3_regs_6_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_1_9 <= stage3_regs_6_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_1_10 <= stage3_regs_6_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_6_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_6_1_11 <= stage3_regs_6_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_7_0_0 <= x_n_30; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_0_1 <= stage3_regs_7_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_0_2 <= stage3_regs_7_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_0_3 <= stage3_regs_7_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_0_4 <= stage3_regs_7_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_0_5 <= stage3_regs_7_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_0_6 <= stage3_regs_7_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_0_7 <= stage3_regs_7_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_0_8 <= stage3_regs_7_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_0_9 <= stage3_regs_7_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_0_10 <= stage3_regs_7_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_0_11 <= stage3_regs_7_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_7_1_0 <= a_2_30; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_1_1 <= stage3_regs_7_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_1_2 <= stage3_regs_7_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_1_3 <= stage3_regs_7_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_1_4 <= stage3_regs_7_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_1_5 <= stage3_regs_7_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_1_6 <= stage3_regs_7_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_1_7 <= stage3_regs_7_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_1_8 <= stage3_regs_7_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_1_9 <= stage3_regs_7_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_1_10 <= stage3_regs_7_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_7_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_7_1_11 <= stage3_regs_7_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_8_0_0 <= x_n_34; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_0_1 <= stage3_regs_8_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_0_2 <= stage3_regs_8_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_0_3 <= stage3_regs_8_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_0_4 <= stage3_regs_8_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_0_5 <= stage3_regs_8_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_0_6 <= stage3_regs_8_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_0_7 <= stage3_regs_8_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_0_8 <= stage3_regs_8_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_0_9 <= stage3_regs_8_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_0_10 <= stage3_regs_8_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_0_11 <= stage3_regs_8_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_8_1_0 <= a_2_34; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_1_1 <= stage3_regs_8_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_1_2 <= stage3_regs_8_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_1_3 <= stage3_regs_8_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_1_4 <= stage3_regs_8_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_1_5 <= stage3_regs_8_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_1_6 <= stage3_regs_8_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_1_7 <= stage3_regs_8_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_1_8 <= stage3_regs_8_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_1_9 <= stage3_regs_8_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_1_10 <= stage3_regs_8_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_8_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_8_1_11 <= stage3_regs_8_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_9_0_0 <= x_n_38; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_0_1 <= stage3_regs_9_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_0_2 <= stage3_regs_9_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_0_3 <= stage3_regs_9_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_0_4 <= stage3_regs_9_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_0_5 <= stage3_regs_9_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_0_6 <= stage3_regs_9_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_0_7 <= stage3_regs_9_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_0_8 <= stage3_regs_9_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_0_9 <= stage3_regs_9_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_0_10 <= stage3_regs_9_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_0_11 <= stage3_regs_9_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_9_1_0 <= a_2_38; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_1_1 <= stage3_regs_9_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_1_2 <= stage3_regs_9_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_1_3 <= stage3_regs_9_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_1_4 <= stage3_regs_9_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_1_5 <= stage3_regs_9_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_1_6 <= stage3_regs_9_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_1_7 <= stage3_regs_9_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_1_8 <= stage3_regs_9_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_1_9 <= stage3_regs_9_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_1_10 <= stage3_regs_9_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_9_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_9_1_11 <= stage3_regs_9_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_10_0_0 <= x_n_42; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_0_1 <= stage3_regs_10_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_0_2 <= stage3_regs_10_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_0_3 <= stage3_regs_10_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_0_4 <= stage3_regs_10_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_0_5 <= stage3_regs_10_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_0_6 <= stage3_regs_10_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_0_7 <= stage3_regs_10_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_0_8 <= stage3_regs_10_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_0_9 <= stage3_regs_10_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_0_10 <= stage3_regs_10_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_0_11 <= stage3_regs_10_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_10_1_0 <= a_2_42; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_1_1 <= stage3_regs_10_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_1_2 <= stage3_regs_10_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_1_3 <= stage3_regs_10_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_1_4 <= stage3_regs_10_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_1_5 <= stage3_regs_10_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_1_6 <= stage3_regs_10_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_1_7 <= stage3_regs_10_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_1_8 <= stage3_regs_10_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_1_9 <= stage3_regs_10_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_1_10 <= stage3_regs_10_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_10_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_10_1_11 <= stage3_regs_10_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_11_0_0 <= x_n_46; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_0_1 <= stage3_regs_11_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_0_2 <= stage3_regs_11_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_0_3 <= stage3_regs_11_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_0_4 <= stage3_regs_11_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_0_5 <= stage3_regs_11_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_0_6 <= stage3_regs_11_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_0_7 <= stage3_regs_11_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_0_8 <= stage3_regs_11_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_0_9 <= stage3_regs_11_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_0_10 <= stage3_regs_11_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_0_11 <= stage3_regs_11_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_11_1_0 <= a_2_46; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_1_1 <= stage3_regs_11_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_1_2 <= stage3_regs_11_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_1_3 <= stage3_regs_11_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_1_4 <= stage3_regs_11_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_1_5 <= stage3_regs_11_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_1_6 <= stage3_regs_11_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_1_7 <= stage3_regs_11_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_1_8 <= stage3_regs_11_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_1_9 <= stage3_regs_11_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_1_10 <= stage3_regs_11_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_11_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_11_1_11 <= stage3_regs_11_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_12_0_0 <= x_n_50; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_0_1 <= stage3_regs_12_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_0_2 <= stage3_regs_12_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_0_3 <= stage3_regs_12_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_0_4 <= stage3_regs_12_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_0_5 <= stage3_regs_12_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_0_6 <= stage3_regs_12_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_0_7 <= stage3_regs_12_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_0_8 <= stage3_regs_12_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_0_9 <= stage3_regs_12_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_0_10 <= stage3_regs_12_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_0_11 <= stage3_regs_12_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_12_1_0 <= a_2_50; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_1_1 <= stage3_regs_12_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_1_2 <= stage3_regs_12_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_1_3 <= stage3_regs_12_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_1_4 <= stage3_regs_12_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_1_5 <= stage3_regs_12_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_1_6 <= stage3_regs_12_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_1_7 <= stage3_regs_12_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_1_8 <= stage3_regs_12_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_1_9 <= stage3_regs_12_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_1_10 <= stage3_regs_12_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_12_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_12_1_11 <= stage3_regs_12_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_13_0_0 <= x_n_54; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_0_1 <= stage3_regs_13_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_0_2 <= stage3_regs_13_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_0_3 <= stage3_regs_13_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_0_4 <= stage3_regs_13_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_0_5 <= stage3_regs_13_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_0_6 <= stage3_regs_13_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_0_7 <= stage3_regs_13_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_0_8 <= stage3_regs_13_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_0_9 <= stage3_regs_13_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_0_10 <= stage3_regs_13_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_0_11 <= stage3_regs_13_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_13_1_0 <= a_2_54; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_1_1 <= stage3_regs_13_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_1_2 <= stage3_regs_13_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_1_3 <= stage3_regs_13_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_1_4 <= stage3_regs_13_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_1_5 <= stage3_regs_13_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_1_6 <= stage3_regs_13_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_1_7 <= stage3_regs_13_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_1_8 <= stage3_regs_13_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_1_9 <= stage3_regs_13_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_1_10 <= stage3_regs_13_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_13_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_13_1_11 <= stage3_regs_13_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_14_0_0 <= x_n_58; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_0_1 <= stage3_regs_14_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_0_2 <= stage3_regs_14_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_0_3 <= stage3_regs_14_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_0_4 <= stage3_regs_14_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_0_5 <= stage3_regs_14_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_0_6 <= stage3_regs_14_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_0_7 <= stage3_regs_14_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_0_8 <= stage3_regs_14_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_0_9 <= stage3_regs_14_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_0_10 <= stage3_regs_14_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_0_11 <= stage3_regs_14_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_14_1_0 <= a_2_58; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_1_1 <= stage3_regs_14_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_1_2 <= stage3_regs_14_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_1_3 <= stage3_regs_14_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_1_4 <= stage3_regs_14_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_1_5 <= stage3_regs_14_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_1_6 <= stage3_regs_14_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_1_7 <= stage3_regs_14_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_1_8 <= stage3_regs_14_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_1_9 <= stage3_regs_14_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_1_10 <= stage3_regs_14_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_14_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_14_1_11 <= stage3_regs_14_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_15_0_0 <= x_n_62; // @[FloatingPointDesigns.scala 2170:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_0_1 <= stage3_regs_15_0_0; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_0_2 <= stage3_regs_15_0_1; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_0_3 <= stage3_regs_15_0_2; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_0_4 <= stage3_regs_15_0_3; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_0_5 <= stage3_regs_15_0_4; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_0_6 <= stage3_regs_15_0_5; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_0_7 <= stage3_regs_15_0_6; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_0_8 <= stage3_regs_15_0_7; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_0_9 <= stage3_regs_15_0_8; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_0_10 <= stage3_regs_15_0_9; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_0_11 <= stage3_regs_15_0_10; // @[FloatingPointDesigns.scala 2123:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2167:26]
      stage3_regs_15_1_0 <= a_2_62; // @[FloatingPointDesigns.scala 2171:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_1_1 <= stage3_regs_15_1_0; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_1_2 <= stage3_regs_15_1_1; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_1_3 <= stage3_regs_15_1_2; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_1_4 <= stage3_regs_15_1_3; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_1_5 <= stage3_regs_15_1_4; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_1_6 <= stage3_regs_15_1_5; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_1_7 <= stage3_regs_15_1_6; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_1_8 <= stage3_regs_15_1_7; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_1_9 <= stage3_regs_15_1_8; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_1_10 <= stage3_regs_15_1_9; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2112:30]
      stage3_regs_15_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2112:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage3_regs_15_1_11 <= stage3_regs_15_1_10; // @[FloatingPointDesigns.scala 2124:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_0_1_0 <= a_2_3; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_0_1_1 <= stage4_regs_0_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_0_1_2 <= stage4_regs_0_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_0_1_3 <= stage4_regs_0_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_0_1_4 <= stage4_regs_0_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_0_1_5 <= stage4_regs_0_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_0_1_6 <= stage4_regs_0_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_0_1_7 <= stage4_regs_0_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_0_1_8 <= stage4_regs_0_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_1_1_0 <= a_2_7; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_1_1_1 <= stage4_regs_1_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_1_1_2 <= stage4_regs_1_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_1_1_3 <= stage4_regs_1_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_1_1_4 <= stage4_regs_1_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_1_1_5 <= stage4_regs_1_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_1_1_6 <= stage4_regs_1_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_1_1_7 <= stage4_regs_1_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_1_1_8 <= stage4_regs_1_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_2_1_0 <= a_2_11; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_2_1_1 <= stage4_regs_2_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_2_1_2 <= stage4_regs_2_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_2_1_3 <= stage4_regs_2_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_2_1_4 <= stage4_regs_2_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_2_1_5 <= stage4_regs_2_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_2_1_6 <= stage4_regs_2_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_2_1_7 <= stage4_regs_2_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_2_1_8 <= stage4_regs_2_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_3_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_3_1_0 <= a_2_15; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_3_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_3_1_1 <= stage4_regs_3_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_3_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_3_1_2 <= stage4_regs_3_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_3_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_3_1_3 <= stage4_regs_3_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_3_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_3_1_4 <= stage4_regs_3_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_3_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_3_1_5 <= stage4_regs_3_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_3_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_3_1_6 <= stage4_regs_3_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_3_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_3_1_7 <= stage4_regs_3_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_3_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_3_1_8 <= stage4_regs_3_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_4_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_4_1_0 <= a_2_19; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_4_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_4_1_1 <= stage4_regs_4_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_4_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_4_1_2 <= stage4_regs_4_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_4_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_4_1_3 <= stage4_regs_4_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_4_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_4_1_4 <= stage4_regs_4_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_4_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_4_1_5 <= stage4_regs_4_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_4_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_4_1_6 <= stage4_regs_4_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_4_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_4_1_7 <= stage4_regs_4_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_4_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_4_1_8 <= stage4_regs_4_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_5_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_5_1_0 <= a_2_23; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_5_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_5_1_1 <= stage4_regs_5_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_5_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_5_1_2 <= stage4_regs_5_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_5_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_5_1_3 <= stage4_regs_5_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_5_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_5_1_4 <= stage4_regs_5_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_5_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_5_1_5 <= stage4_regs_5_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_5_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_5_1_6 <= stage4_regs_5_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_5_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_5_1_7 <= stage4_regs_5_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_5_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_5_1_8 <= stage4_regs_5_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_6_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_6_1_0 <= a_2_27; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_6_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_6_1_1 <= stage4_regs_6_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_6_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_6_1_2 <= stage4_regs_6_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_6_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_6_1_3 <= stage4_regs_6_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_6_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_6_1_4 <= stage4_regs_6_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_6_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_6_1_5 <= stage4_regs_6_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_6_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_6_1_6 <= stage4_regs_6_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_6_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_6_1_7 <= stage4_regs_6_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_6_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_6_1_8 <= stage4_regs_6_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_7_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_7_1_0 <= a_2_31; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_7_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_7_1_1 <= stage4_regs_7_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_7_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_7_1_2 <= stage4_regs_7_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_7_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_7_1_3 <= stage4_regs_7_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_7_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_7_1_4 <= stage4_regs_7_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_7_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_7_1_5 <= stage4_regs_7_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_7_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_7_1_6 <= stage4_regs_7_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_7_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_7_1_7 <= stage4_regs_7_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_7_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_7_1_8 <= stage4_regs_7_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_8_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_8_1_0 <= a_2_35; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_8_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_8_1_1 <= stage4_regs_8_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_8_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_8_1_2 <= stage4_regs_8_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_8_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_8_1_3 <= stage4_regs_8_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_8_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_8_1_4 <= stage4_regs_8_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_8_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_8_1_5 <= stage4_regs_8_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_8_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_8_1_6 <= stage4_regs_8_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_8_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_8_1_7 <= stage4_regs_8_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_8_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_8_1_8 <= stage4_regs_8_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_9_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_9_1_0 <= a_2_39; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_9_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_9_1_1 <= stage4_regs_9_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_9_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_9_1_2 <= stage4_regs_9_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_9_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_9_1_3 <= stage4_regs_9_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_9_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_9_1_4 <= stage4_regs_9_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_9_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_9_1_5 <= stage4_regs_9_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_9_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_9_1_6 <= stage4_regs_9_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_9_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_9_1_7 <= stage4_regs_9_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_9_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_9_1_8 <= stage4_regs_9_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_10_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_10_1_0 <= a_2_43; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_10_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_10_1_1 <= stage4_regs_10_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_10_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_10_1_2 <= stage4_regs_10_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_10_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_10_1_3 <= stage4_regs_10_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_10_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_10_1_4 <= stage4_regs_10_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_10_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_10_1_5 <= stage4_regs_10_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_10_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_10_1_6 <= stage4_regs_10_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_10_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_10_1_7 <= stage4_regs_10_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_10_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_10_1_8 <= stage4_regs_10_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_11_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_11_1_0 <= a_2_47; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_11_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_11_1_1 <= stage4_regs_11_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_11_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_11_1_2 <= stage4_regs_11_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_11_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_11_1_3 <= stage4_regs_11_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_11_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_11_1_4 <= stage4_regs_11_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_11_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_11_1_5 <= stage4_regs_11_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_11_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_11_1_6 <= stage4_regs_11_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_11_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_11_1_7 <= stage4_regs_11_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_11_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_11_1_8 <= stage4_regs_11_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_12_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_12_1_0 <= a_2_51; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_12_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_12_1_1 <= stage4_regs_12_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_12_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_12_1_2 <= stage4_regs_12_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_12_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_12_1_3 <= stage4_regs_12_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_12_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_12_1_4 <= stage4_regs_12_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_12_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_12_1_5 <= stage4_regs_12_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_12_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_12_1_6 <= stage4_regs_12_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_12_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_12_1_7 <= stage4_regs_12_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_12_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_12_1_8 <= stage4_regs_12_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_13_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_13_1_0 <= a_2_55; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_13_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_13_1_1 <= stage4_regs_13_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_13_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_13_1_2 <= stage4_regs_13_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_13_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_13_1_3 <= stage4_regs_13_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_13_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_13_1_4 <= stage4_regs_13_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_13_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_13_1_5 <= stage4_regs_13_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_13_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_13_1_6 <= stage4_regs_13_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_13_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_13_1_7 <= stage4_regs_13_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_13_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_13_1_8 <= stage4_regs_13_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_14_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_14_1_0 <= a_2_59; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_14_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_14_1_1 <= stage4_regs_14_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_14_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_14_1_2 <= stage4_regs_14_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_14_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_14_1_3 <= stage4_regs_14_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_14_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_14_1_4 <= stage4_regs_14_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_14_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_14_1_5 <= stage4_regs_14_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_14_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_14_1_6 <= stage4_regs_14_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_14_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_14_1_7 <= stage4_regs_14_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_14_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_14_1_8 <= stage4_regs_14_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_15_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2176:26]
      stage4_regs_15_1_0 <= a_2_63; // @[FloatingPointDesigns.scala 2178:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_15_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_15_1_1 <= stage4_regs_15_1_0; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_15_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_15_1_2 <= stage4_regs_15_1_1; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_15_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_15_1_3 <= stage4_regs_15_1_2; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_15_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_15_1_4 <= stage4_regs_15_1_3; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_15_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_15_1_5 <= stage4_regs_15_1_4; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_15_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_15_1_6 <= stage4_regs_15_1_5; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_15_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_15_1_7 <= stage4_regs_15_1_6; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2113:30]
      stage4_regs_15_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2113:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2121:22]
      stage4_regs_15_1_8 <= stage4_regs_15_1_7; // @[FloatingPointDesigns.scala 2130:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2184:31]
      a_2_isr_to_r <= 32'h0; // @[FloatingPointDesigns.scala 2184:31]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2186:20]
      a_2_isr_to_r <= _a_2_isr_to_r_T_6; // @[FloatingPointDesigns.scala 2187:20]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2185:34]
      transition_regs_0 <= 32'h0; // @[FloatingPointDesigns.scala 2185:34]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2186:20]
      transition_regs_0 <= a_2_isr_to_r; // @[FloatingPointDesigns.scala 2188:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2185:34]
      transition_regs_1 <= 32'h0; // @[FloatingPointDesigns.scala 2185:34]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2186:20]
      transition_regs_1 <= transition_regs_0; // @[FloatingPointDesigns.scala 2190:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2185:34]
      transition_regs_2 <= 32'h0; // @[FloatingPointDesigns.scala 2185:34]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2186:20]
      transition_regs_2 <= transition_regs_1; // @[FloatingPointDesigns.scala 2190:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2185:34]
      transition_regs_3 <= 32'h0; // @[FloatingPointDesigns.scala 2185:34]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2186:20]
      transition_regs_3 <= transition_regs_2; // @[FloatingPointDesigns.scala 2190:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2185:34]
      transition_regs_4 <= 32'h0; // @[FloatingPointDesigns.scala 2185:34]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2186:20]
      transition_regs_4 <= transition_regs_3; // @[FloatingPointDesigns.scala 2190:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2185:34]
      transition_regs_5 <= 32'h0; // @[FloatingPointDesigns.scala 2185:34]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2186:20]
      transition_regs_5 <= transition_regs_4; // @[FloatingPointDesigns.scala 2190:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2185:34]
      transition_regs_6 <= 32'h0; // @[FloatingPointDesigns.scala 2185:34]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2186:20]
      transition_regs_6 <= transition_regs_5; // @[FloatingPointDesigns.scala 2190:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2185:34]
      transition_regs_7 <= 32'h0; // @[FloatingPointDesigns.scala 2185:34]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2186:20]
      transition_regs_7 <= transition_regs_6; // @[FloatingPointDesigns.scala 2190:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2185:34]
      transition_regs_8 <= 32'h0; // @[FloatingPointDesigns.scala 2185:34]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2186:20]
      transition_regs_8 <= transition_regs_7; // @[FloatingPointDesigns.scala 2190:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_0 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2226:28]
      x_n_r_0 <= multiplier4_io_out_s; // @[FloatingPointDesigns.scala 2227:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_1 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_1 <= stage1_regs_r_0_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_3 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_3 <= FP_multiplier_10ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_4 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_4 <= stage1_regs_r_1_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_6 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_6 <= FP_multiplier_10ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_7 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_7 <= stage1_regs_r_2_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_9 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_9 <= FP_multiplier_10ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_10 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_10 <= stage1_regs_r_3_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_12 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_12 <= FP_multiplier_10ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_13 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_13 <= stage1_regs_r_4_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_15 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_15 <= FP_multiplier_10ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_16 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_16 <= stage1_regs_r_5_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_18 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_18 <= FP_multiplier_10ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_19 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_19 <= stage1_regs_r_6_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_21 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_21 <= FP_multiplier_10ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_22 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_22 <= stage1_regs_r_7_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_24 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_24 <= FP_multiplier_10ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_25 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_25 <= stage1_regs_r_8_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_27 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_27 <= FP_multiplier_10ccs_65_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_28 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_28 <= stage1_regs_r_9_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_30 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_30 <= FP_multiplier_10ccs_67_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_31 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_31 <= stage1_regs_r_10_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_33 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_33 <= FP_multiplier_10ccs_69_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_34 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_34 <= stage1_regs_r_11_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_36 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_36 <= FP_multiplier_10ccs_71_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_37 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_37 <= stage1_regs_r_12_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_39 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_39 <= FP_multiplier_10ccs_73_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_40 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_40 <= stage1_regs_r_13_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_42 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_42 <= FP_multiplier_10ccs_75_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_43 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_43 <= stage1_regs_r_14_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_45 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_45 <= FP_multiplier_10ccs_77_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_46 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_46 <= stage1_regs_r_15_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_48 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      x_n_r_48 <= FP_multiplier_10ccs_79_io_out_s; // @[FloatingPointDesigns.scala 2236:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2201:24]
      x_n_r_49 <= 32'h0; // @[FloatingPointDesigns.scala 2201:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      x_n_r_49 <= stage1_regs_r_16_0_8; // @[FloatingPointDesigns.scala 2249:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_0 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2226:28]
      a_2_r_0 <= transition_regs_8; // @[FloatingPointDesigns.scala 2228:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_1 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_1 <= stage1_regs_r_0_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_2 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_2 <= stage2_regs_r_0_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_3 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_3 <= stage3_regs_r_0_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_4 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_4 <= stage1_regs_r_1_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_5 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_5 <= stage2_regs_r_1_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_6 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_6 <= stage3_regs_r_1_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_7 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_7 <= stage1_regs_r_2_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_8 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_8 <= stage2_regs_r_2_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_9 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_9 <= stage3_regs_r_2_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_10 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_10 <= stage1_regs_r_3_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_11 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_11 <= stage2_regs_r_3_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_12 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_12 <= stage3_regs_r_3_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_13 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_13 <= stage1_regs_r_4_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_14 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_14 <= stage2_regs_r_4_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_15 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_15 <= stage3_regs_r_4_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_16 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_16 <= stage1_regs_r_5_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_17 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_17 <= stage2_regs_r_5_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_18 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_18 <= stage3_regs_r_5_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_19 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_19 <= stage1_regs_r_6_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_20 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_20 <= stage2_regs_r_6_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_21 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_21 <= stage3_regs_r_6_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_22 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_22 <= stage1_regs_r_7_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_23 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_23 <= stage2_regs_r_7_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_24 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_24 <= stage3_regs_r_7_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_25 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_25 <= stage1_regs_r_8_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_26 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_26 <= stage2_regs_r_8_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_27 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_27 <= stage3_regs_r_8_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_28 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_28 <= stage1_regs_r_9_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_29 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_29 <= stage2_regs_r_9_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_30 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_30 <= stage3_regs_r_9_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_31 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_31 <= stage1_regs_r_10_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_32 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_32 <= stage2_regs_r_10_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_33 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_33 <= stage3_regs_r_10_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_34 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_34 <= stage1_regs_r_11_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_35 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_35 <= stage2_regs_r_11_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_36 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_36 <= stage3_regs_r_11_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_37 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_37 <= stage1_regs_r_12_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_38 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_38 <= stage2_regs_r_12_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_39 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_39 <= stage3_regs_r_12_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_40 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_40 <= stage1_regs_r_13_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_41 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_41 <= stage2_regs_r_13_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_42 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_42 <= stage3_regs_r_13_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_43 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_43 <= stage1_regs_r_14_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_44 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_44 <= stage2_regs_r_14_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_45 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_45 <= stage3_regs_r_14_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_46 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_46 <= stage1_regs_r_15_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_47 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_47 <= stage2_regs_r_15_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_48 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      a_2_r_48 <= stage3_regs_r_15_1_8; // @[FloatingPointDesigns.scala 2237:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_49 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      a_2_r_49 <= stage1_regs_r_16_1_8; // @[FloatingPointDesigns.scala 2248:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2202:24]
      a_2_r_50 <= 32'h0; // @[FloatingPointDesigns.scala 2202:24]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      a_2_r_50 <= stage2_regs_r_16_1_11; // @[FloatingPointDesigns.scala 2257:30]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2226:28]
      stage1_regs_r_0_0_0 <= x_n_r_0; // @[FloatingPointDesigns.scala 2229:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_0_1 <= stage1_regs_r_0_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_0_2 <= stage1_regs_r_0_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_0_3 <= stage1_regs_r_0_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_0_4 <= stage1_regs_r_0_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_0_5 <= stage1_regs_r_0_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_0_6 <= stage1_regs_r_0_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_0_7 <= stage1_regs_r_0_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_0_8 <= stage1_regs_r_0_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2226:28]
      stage1_regs_r_0_1_0 <= a_2_r_0; // @[FloatingPointDesigns.scala 2230:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_1_1 <= stage1_regs_r_0_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_1_2 <= stage1_regs_r_0_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_1_3 <= stage1_regs_r_0_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_1_4 <= stage1_regs_r_0_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_1_5 <= stage1_regs_r_0_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_1_6 <= stage1_regs_r_0_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_1_7 <= stage1_regs_r_0_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_0_1_8 <= stage1_regs_r_0_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_1_0_0 <= x_n_r_3; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_0_1 <= stage1_regs_r_1_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_0_2 <= stage1_regs_r_1_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_0_3 <= stage1_regs_r_1_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_0_4 <= stage1_regs_r_1_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_0_5 <= stage1_regs_r_1_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_0_6 <= stage1_regs_r_1_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_0_7 <= stage1_regs_r_1_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_0_8 <= stage1_regs_r_1_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_1_1_0 <= a_2_r_3; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_1_1 <= stage1_regs_r_1_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_1_2 <= stage1_regs_r_1_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_1_3 <= stage1_regs_r_1_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_1_4 <= stage1_regs_r_1_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_1_5 <= stage1_regs_r_1_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_1_6 <= stage1_regs_r_1_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_1_7 <= stage1_regs_r_1_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_1_1_8 <= stage1_regs_r_1_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_2_0_0 <= x_n_r_6; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_0_1 <= stage1_regs_r_2_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_0_2 <= stage1_regs_r_2_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_0_3 <= stage1_regs_r_2_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_0_4 <= stage1_regs_r_2_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_0_5 <= stage1_regs_r_2_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_0_6 <= stage1_regs_r_2_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_0_7 <= stage1_regs_r_2_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_0_8 <= stage1_regs_r_2_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_2_1_0 <= a_2_r_6; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_1_1 <= stage1_regs_r_2_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_1_2 <= stage1_regs_r_2_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_1_3 <= stage1_regs_r_2_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_1_4 <= stage1_regs_r_2_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_1_5 <= stage1_regs_r_2_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_1_6 <= stage1_regs_r_2_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_1_7 <= stage1_regs_r_2_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_2_1_8 <= stage1_regs_r_2_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_3_0_0 <= x_n_r_9; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_0_1 <= stage1_regs_r_3_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_0_2 <= stage1_regs_r_3_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_0_3 <= stage1_regs_r_3_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_0_4 <= stage1_regs_r_3_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_0_5 <= stage1_regs_r_3_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_0_6 <= stage1_regs_r_3_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_0_7 <= stage1_regs_r_3_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_0_8 <= stage1_regs_r_3_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_3_1_0 <= a_2_r_9; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_1_1 <= stage1_regs_r_3_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_1_2 <= stage1_regs_r_3_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_1_3 <= stage1_regs_r_3_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_1_4 <= stage1_regs_r_3_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_1_5 <= stage1_regs_r_3_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_1_6 <= stage1_regs_r_3_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_1_7 <= stage1_regs_r_3_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_3_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_3_1_8 <= stage1_regs_r_3_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_4_0_0 <= x_n_r_12; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_0_1 <= stage1_regs_r_4_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_0_2 <= stage1_regs_r_4_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_0_3 <= stage1_regs_r_4_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_0_4 <= stage1_regs_r_4_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_0_5 <= stage1_regs_r_4_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_0_6 <= stage1_regs_r_4_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_0_7 <= stage1_regs_r_4_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_0_8 <= stage1_regs_r_4_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_4_1_0 <= a_2_r_12; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_1_1 <= stage1_regs_r_4_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_1_2 <= stage1_regs_r_4_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_1_3 <= stage1_regs_r_4_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_1_4 <= stage1_regs_r_4_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_1_5 <= stage1_regs_r_4_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_1_6 <= stage1_regs_r_4_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_1_7 <= stage1_regs_r_4_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_4_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_4_1_8 <= stage1_regs_r_4_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_5_0_0 <= x_n_r_15; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_0_1 <= stage1_regs_r_5_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_0_2 <= stage1_regs_r_5_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_0_3 <= stage1_regs_r_5_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_0_4 <= stage1_regs_r_5_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_0_5 <= stage1_regs_r_5_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_0_6 <= stage1_regs_r_5_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_0_7 <= stage1_regs_r_5_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_0_8 <= stage1_regs_r_5_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_5_1_0 <= a_2_r_15; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_1_1 <= stage1_regs_r_5_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_1_2 <= stage1_regs_r_5_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_1_3 <= stage1_regs_r_5_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_1_4 <= stage1_regs_r_5_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_1_5 <= stage1_regs_r_5_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_1_6 <= stage1_regs_r_5_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_1_7 <= stage1_regs_r_5_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_5_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_5_1_8 <= stage1_regs_r_5_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_6_0_0 <= x_n_r_18; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_0_1 <= stage1_regs_r_6_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_0_2 <= stage1_regs_r_6_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_0_3 <= stage1_regs_r_6_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_0_4 <= stage1_regs_r_6_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_0_5 <= stage1_regs_r_6_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_0_6 <= stage1_regs_r_6_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_0_7 <= stage1_regs_r_6_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_0_8 <= stage1_regs_r_6_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_6_1_0 <= a_2_r_18; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_1_1 <= stage1_regs_r_6_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_1_2 <= stage1_regs_r_6_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_1_3 <= stage1_regs_r_6_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_1_4 <= stage1_regs_r_6_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_1_5 <= stage1_regs_r_6_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_1_6 <= stage1_regs_r_6_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_1_7 <= stage1_regs_r_6_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_6_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_6_1_8 <= stage1_regs_r_6_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_7_0_0 <= x_n_r_21; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_0_1 <= stage1_regs_r_7_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_0_2 <= stage1_regs_r_7_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_0_3 <= stage1_regs_r_7_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_0_4 <= stage1_regs_r_7_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_0_5 <= stage1_regs_r_7_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_0_6 <= stage1_regs_r_7_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_0_7 <= stage1_regs_r_7_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_0_8 <= stage1_regs_r_7_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_7_1_0 <= a_2_r_21; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_1_1 <= stage1_regs_r_7_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_1_2 <= stage1_regs_r_7_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_1_3 <= stage1_regs_r_7_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_1_4 <= stage1_regs_r_7_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_1_5 <= stage1_regs_r_7_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_1_6 <= stage1_regs_r_7_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_1_7 <= stage1_regs_r_7_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_7_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_7_1_8 <= stage1_regs_r_7_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_8_0_0 <= x_n_r_24; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_0_1 <= stage1_regs_r_8_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_0_2 <= stage1_regs_r_8_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_0_3 <= stage1_regs_r_8_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_0_4 <= stage1_regs_r_8_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_0_5 <= stage1_regs_r_8_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_0_6 <= stage1_regs_r_8_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_0_7 <= stage1_regs_r_8_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_0_8 <= stage1_regs_r_8_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_8_1_0 <= a_2_r_24; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_1_1 <= stage1_regs_r_8_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_1_2 <= stage1_regs_r_8_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_1_3 <= stage1_regs_r_8_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_1_4 <= stage1_regs_r_8_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_1_5 <= stage1_regs_r_8_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_1_6 <= stage1_regs_r_8_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_1_7 <= stage1_regs_r_8_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_8_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_8_1_8 <= stage1_regs_r_8_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_9_0_0 <= x_n_r_27; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_0_1 <= stage1_regs_r_9_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_0_2 <= stage1_regs_r_9_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_0_3 <= stage1_regs_r_9_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_0_4 <= stage1_regs_r_9_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_0_5 <= stage1_regs_r_9_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_0_6 <= stage1_regs_r_9_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_0_7 <= stage1_regs_r_9_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_0_8 <= stage1_regs_r_9_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_9_1_0 <= a_2_r_27; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_1_1 <= stage1_regs_r_9_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_1_2 <= stage1_regs_r_9_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_1_3 <= stage1_regs_r_9_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_1_4 <= stage1_regs_r_9_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_1_5 <= stage1_regs_r_9_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_1_6 <= stage1_regs_r_9_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_1_7 <= stage1_regs_r_9_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_9_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_9_1_8 <= stage1_regs_r_9_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_10_0_0 <= x_n_r_30; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_0_1 <= stage1_regs_r_10_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_0_2 <= stage1_regs_r_10_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_0_3 <= stage1_regs_r_10_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_0_4 <= stage1_regs_r_10_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_0_5 <= stage1_regs_r_10_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_0_6 <= stage1_regs_r_10_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_0_7 <= stage1_regs_r_10_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_0_8 <= stage1_regs_r_10_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_10_1_0 <= a_2_r_30; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_1_1 <= stage1_regs_r_10_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_1_2 <= stage1_regs_r_10_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_1_3 <= stage1_regs_r_10_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_1_4 <= stage1_regs_r_10_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_1_5 <= stage1_regs_r_10_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_1_6 <= stage1_regs_r_10_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_1_7 <= stage1_regs_r_10_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_10_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_10_1_8 <= stage1_regs_r_10_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_11_0_0 <= x_n_r_33; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_0_1 <= stage1_regs_r_11_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_0_2 <= stage1_regs_r_11_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_0_3 <= stage1_regs_r_11_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_0_4 <= stage1_regs_r_11_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_0_5 <= stage1_regs_r_11_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_0_6 <= stage1_regs_r_11_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_0_7 <= stage1_regs_r_11_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_0_8 <= stage1_regs_r_11_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_11_1_0 <= a_2_r_33; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_1_1 <= stage1_regs_r_11_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_1_2 <= stage1_regs_r_11_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_1_3 <= stage1_regs_r_11_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_1_4 <= stage1_regs_r_11_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_1_5 <= stage1_regs_r_11_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_1_6 <= stage1_regs_r_11_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_1_7 <= stage1_regs_r_11_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_11_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_11_1_8 <= stage1_regs_r_11_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_12_0_0 <= x_n_r_36; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_0_1 <= stage1_regs_r_12_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_0_2 <= stage1_regs_r_12_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_0_3 <= stage1_regs_r_12_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_0_4 <= stage1_regs_r_12_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_0_5 <= stage1_regs_r_12_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_0_6 <= stage1_regs_r_12_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_0_7 <= stage1_regs_r_12_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_0_8 <= stage1_regs_r_12_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_12_1_0 <= a_2_r_36; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_1_1 <= stage1_regs_r_12_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_1_2 <= stage1_regs_r_12_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_1_3 <= stage1_regs_r_12_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_1_4 <= stage1_regs_r_12_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_1_5 <= stage1_regs_r_12_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_1_6 <= stage1_regs_r_12_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_1_7 <= stage1_regs_r_12_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_12_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_12_1_8 <= stage1_regs_r_12_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_13_0_0 <= x_n_r_39; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_0_1 <= stage1_regs_r_13_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_0_2 <= stage1_regs_r_13_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_0_3 <= stage1_regs_r_13_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_0_4 <= stage1_regs_r_13_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_0_5 <= stage1_regs_r_13_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_0_6 <= stage1_regs_r_13_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_0_7 <= stage1_regs_r_13_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_0_8 <= stage1_regs_r_13_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_13_1_0 <= a_2_r_39; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_1_1 <= stage1_regs_r_13_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_1_2 <= stage1_regs_r_13_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_1_3 <= stage1_regs_r_13_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_1_4 <= stage1_regs_r_13_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_1_5 <= stage1_regs_r_13_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_1_6 <= stage1_regs_r_13_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_1_7 <= stage1_regs_r_13_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_13_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_13_1_8 <= stage1_regs_r_13_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_14_0_0 <= x_n_r_42; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_0_1 <= stage1_regs_r_14_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_0_2 <= stage1_regs_r_14_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_0_3 <= stage1_regs_r_14_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_0_4 <= stage1_regs_r_14_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_0_5 <= stage1_regs_r_14_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_0_6 <= stage1_regs_r_14_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_0_7 <= stage1_regs_r_14_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_0_8 <= stage1_regs_r_14_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_14_1_0 <= a_2_r_42; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_1_1 <= stage1_regs_r_14_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_1_2 <= stage1_regs_r_14_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_1_3 <= stage1_regs_r_14_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_1_4 <= stage1_regs_r_14_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_1_5 <= stage1_regs_r_14_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_1_6 <= stage1_regs_r_14_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_1_7 <= stage1_regs_r_14_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_14_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_14_1_8 <= stage1_regs_r_14_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_15_0_0 <= x_n_r_45; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_0_1 <= stage1_regs_r_15_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_0_2 <= stage1_regs_r_15_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_0_3 <= stage1_regs_r_15_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_0_4 <= stage1_regs_r_15_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_0_5 <= stage1_regs_r_15_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_0_6 <= stage1_regs_r_15_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_0_7 <= stage1_regs_r_15_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_0_8 <= stage1_regs_r_15_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_15_1_0 <= a_2_r_45; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_1_1 <= stage1_regs_r_15_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_1_2 <= stage1_regs_r_15_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_1_3 <= stage1_regs_r_15_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_1_4 <= stage1_regs_r_15_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_1_5 <= stage1_regs_r_15_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_1_6 <= stage1_regs_r_15_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_1_7 <= stage1_regs_r_15_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_15_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_15_1_8 <= stage1_regs_r_15_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_16_0_0 <= x_n_r_48; // @[FloatingPointDesigns.scala 2238:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_0_1 <= stage1_regs_r_16_0_0; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_0_2 <= stage1_regs_r_16_0_1; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_0_3 <= stage1_regs_r_16_0_2; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_0_4 <= stage1_regs_r_16_0_3; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_0_5 <= stage1_regs_r_16_0_4; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_0_6 <= stage1_regs_r_16_0_5; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_0_7 <= stage1_regs_r_16_0_6; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_0_8 <= stage1_regs_r_16_0_7; // @[FloatingPointDesigns.scala 2217:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2235:28]
      stage1_regs_r_16_1_0 <= a_2_r_48; // @[FloatingPointDesigns.scala 2239:38]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_1_1 <= stage1_regs_r_16_1_0; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_1_2 <= stage1_regs_r_16_1_1; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_1_3 <= stage1_regs_r_16_1_2; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_1_4 <= stage1_regs_r_16_1_3; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_1_5 <= stage1_regs_r_16_1_4; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_1_6 <= stage1_regs_r_16_1_5; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_1_7 <= stage1_regs_r_16_1_6; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2203:32]
      stage1_regs_r_16_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2203:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage1_regs_r_16_1_8 <= stage1_regs_r_16_1_7; // @[FloatingPointDesigns.scala 2218:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_0_0_0 <= x_n_r_1; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_0_1 <= stage2_regs_r_0_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_0_2 <= stage2_regs_r_0_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_0_3 <= stage2_regs_r_0_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_0_4 <= stage2_regs_r_0_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_0_5 <= stage2_regs_r_0_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_0_6 <= stage2_regs_r_0_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_0_7 <= stage2_regs_r_0_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_0_8 <= stage2_regs_r_0_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_0_9 <= stage2_regs_r_0_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_0_10 <= stage2_regs_r_0_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_0_11 <= stage2_regs_r_0_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_0_1_0 <= a_2_r_1; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_1_1 <= stage2_regs_r_0_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_1_2 <= stage2_regs_r_0_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_1_3 <= stage2_regs_r_0_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_1_4 <= stage2_regs_r_0_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_1_5 <= stage2_regs_r_0_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_1_6 <= stage2_regs_r_0_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_1_7 <= stage2_regs_r_0_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_1_8 <= stage2_regs_r_0_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_1_9 <= stage2_regs_r_0_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_1_10 <= stage2_regs_r_0_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_0_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_0_1_11 <= stage2_regs_r_0_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_1_0_0 <= x_n_r_4; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_0_1 <= stage2_regs_r_1_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_0_2 <= stage2_regs_r_1_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_0_3 <= stage2_regs_r_1_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_0_4 <= stage2_regs_r_1_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_0_5 <= stage2_regs_r_1_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_0_6 <= stage2_regs_r_1_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_0_7 <= stage2_regs_r_1_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_0_8 <= stage2_regs_r_1_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_0_9 <= stage2_regs_r_1_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_0_10 <= stage2_regs_r_1_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_0_11 <= stage2_regs_r_1_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_1_1_0 <= a_2_r_4; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_1_1 <= stage2_regs_r_1_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_1_2 <= stage2_regs_r_1_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_1_3 <= stage2_regs_r_1_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_1_4 <= stage2_regs_r_1_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_1_5 <= stage2_regs_r_1_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_1_6 <= stage2_regs_r_1_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_1_7 <= stage2_regs_r_1_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_1_8 <= stage2_regs_r_1_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_1_9 <= stage2_regs_r_1_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_1_10 <= stage2_regs_r_1_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_1_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_1_1_11 <= stage2_regs_r_1_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_2_0_0 <= x_n_r_7; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_0_1 <= stage2_regs_r_2_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_0_2 <= stage2_regs_r_2_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_0_3 <= stage2_regs_r_2_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_0_4 <= stage2_regs_r_2_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_0_5 <= stage2_regs_r_2_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_0_6 <= stage2_regs_r_2_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_0_7 <= stage2_regs_r_2_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_0_8 <= stage2_regs_r_2_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_0_9 <= stage2_regs_r_2_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_0_10 <= stage2_regs_r_2_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_0_11 <= stage2_regs_r_2_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_2_1_0 <= a_2_r_7; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_1_1 <= stage2_regs_r_2_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_1_2 <= stage2_regs_r_2_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_1_3 <= stage2_regs_r_2_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_1_4 <= stage2_regs_r_2_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_1_5 <= stage2_regs_r_2_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_1_6 <= stage2_regs_r_2_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_1_7 <= stage2_regs_r_2_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_1_8 <= stage2_regs_r_2_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_1_9 <= stage2_regs_r_2_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_1_10 <= stage2_regs_r_2_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_2_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_2_1_11 <= stage2_regs_r_2_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_3_0_0 <= x_n_r_10; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_0_1 <= stage2_regs_r_3_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_0_2 <= stage2_regs_r_3_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_0_3 <= stage2_regs_r_3_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_0_4 <= stage2_regs_r_3_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_0_5 <= stage2_regs_r_3_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_0_6 <= stage2_regs_r_3_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_0_7 <= stage2_regs_r_3_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_0_8 <= stage2_regs_r_3_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_0_9 <= stage2_regs_r_3_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_0_10 <= stage2_regs_r_3_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_0_11 <= stage2_regs_r_3_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_3_1_0 <= a_2_r_10; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_1_1 <= stage2_regs_r_3_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_1_2 <= stage2_regs_r_3_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_1_3 <= stage2_regs_r_3_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_1_4 <= stage2_regs_r_3_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_1_5 <= stage2_regs_r_3_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_1_6 <= stage2_regs_r_3_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_1_7 <= stage2_regs_r_3_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_1_8 <= stage2_regs_r_3_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_1_9 <= stage2_regs_r_3_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_1_10 <= stage2_regs_r_3_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_3_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_3_1_11 <= stage2_regs_r_3_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_4_0_0 <= x_n_r_13; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_0_1 <= stage2_regs_r_4_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_0_2 <= stage2_regs_r_4_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_0_3 <= stage2_regs_r_4_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_0_4 <= stage2_regs_r_4_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_0_5 <= stage2_regs_r_4_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_0_6 <= stage2_regs_r_4_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_0_7 <= stage2_regs_r_4_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_0_8 <= stage2_regs_r_4_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_0_9 <= stage2_regs_r_4_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_0_10 <= stage2_regs_r_4_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_0_11 <= stage2_regs_r_4_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_4_1_0 <= a_2_r_13; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_1_1 <= stage2_regs_r_4_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_1_2 <= stage2_regs_r_4_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_1_3 <= stage2_regs_r_4_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_1_4 <= stage2_regs_r_4_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_1_5 <= stage2_regs_r_4_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_1_6 <= stage2_regs_r_4_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_1_7 <= stage2_regs_r_4_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_1_8 <= stage2_regs_r_4_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_1_9 <= stage2_regs_r_4_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_1_10 <= stage2_regs_r_4_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_4_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_4_1_11 <= stage2_regs_r_4_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_5_0_0 <= x_n_r_16; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_0_1 <= stage2_regs_r_5_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_0_2 <= stage2_regs_r_5_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_0_3 <= stage2_regs_r_5_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_0_4 <= stage2_regs_r_5_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_0_5 <= stage2_regs_r_5_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_0_6 <= stage2_regs_r_5_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_0_7 <= stage2_regs_r_5_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_0_8 <= stage2_regs_r_5_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_0_9 <= stage2_regs_r_5_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_0_10 <= stage2_regs_r_5_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_0_11 <= stage2_regs_r_5_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_5_1_0 <= a_2_r_16; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_1_1 <= stage2_regs_r_5_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_1_2 <= stage2_regs_r_5_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_1_3 <= stage2_regs_r_5_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_1_4 <= stage2_regs_r_5_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_1_5 <= stage2_regs_r_5_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_1_6 <= stage2_regs_r_5_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_1_7 <= stage2_regs_r_5_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_1_8 <= stage2_regs_r_5_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_1_9 <= stage2_regs_r_5_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_1_10 <= stage2_regs_r_5_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_5_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_5_1_11 <= stage2_regs_r_5_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_6_0_0 <= x_n_r_19; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_0_1 <= stage2_regs_r_6_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_0_2 <= stage2_regs_r_6_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_0_3 <= stage2_regs_r_6_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_0_4 <= stage2_regs_r_6_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_0_5 <= stage2_regs_r_6_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_0_6 <= stage2_regs_r_6_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_0_7 <= stage2_regs_r_6_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_0_8 <= stage2_regs_r_6_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_0_9 <= stage2_regs_r_6_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_0_10 <= stage2_regs_r_6_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_0_11 <= stage2_regs_r_6_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_6_1_0 <= a_2_r_19; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_1_1 <= stage2_regs_r_6_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_1_2 <= stage2_regs_r_6_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_1_3 <= stage2_regs_r_6_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_1_4 <= stage2_regs_r_6_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_1_5 <= stage2_regs_r_6_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_1_6 <= stage2_regs_r_6_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_1_7 <= stage2_regs_r_6_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_1_8 <= stage2_regs_r_6_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_1_9 <= stage2_regs_r_6_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_1_10 <= stage2_regs_r_6_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_6_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_6_1_11 <= stage2_regs_r_6_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_7_0_0 <= x_n_r_22; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_0_1 <= stage2_regs_r_7_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_0_2 <= stage2_regs_r_7_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_0_3 <= stage2_regs_r_7_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_0_4 <= stage2_regs_r_7_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_0_5 <= stage2_regs_r_7_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_0_6 <= stage2_regs_r_7_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_0_7 <= stage2_regs_r_7_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_0_8 <= stage2_regs_r_7_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_0_9 <= stage2_regs_r_7_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_0_10 <= stage2_regs_r_7_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_0_11 <= stage2_regs_r_7_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_7_1_0 <= a_2_r_22; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_1_1 <= stage2_regs_r_7_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_1_2 <= stage2_regs_r_7_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_1_3 <= stage2_regs_r_7_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_1_4 <= stage2_regs_r_7_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_1_5 <= stage2_regs_r_7_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_1_6 <= stage2_regs_r_7_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_1_7 <= stage2_regs_r_7_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_1_8 <= stage2_regs_r_7_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_1_9 <= stage2_regs_r_7_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_1_10 <= stage2_regs_r_7_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_7_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_7_1_11 <= stage2_regs_r_7_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_8_0_0 <= x_n_r_25; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_0_1 <= stage2_regs_r_8_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_0_2 <= stage2_regs_r_8_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_0_3 <= stage2_regs_r_8_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_0_4 <= stage2_regs_r_8_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_0_5 <= stage2_regs_r_8_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_0_6 <= stage2_regs_r_8_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_0_7 <= stage2_regs_r_8_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_0_8 <= stage2_regs_r_8_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_0_9 <= stage2_regs_r_8_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_0_10 <= stage2_regs_r_8_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_0_11 <= stage2_regs_r_8_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_8_1_0 <= a_2_r_25; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_1_1 <= stage2_regs_r_8_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_1_2 <= stage2_regs_r_8_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_1_3 <= stage2_regs_r_8_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_1_4 <= stage2_regs_r_8_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_1_5 <= stage2_regs_r_8_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_1_6 <= stage2_regs_r_8_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_1_7 <= stage2_regs_r_8_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_1_8 <= stage2_regs_r_8_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_1_9 <= stage2_regs_r_8_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_1_10 <= stage2_regs_r_8_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_8_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_8_1_11 <= stage2_regs_r_8_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_9_0_0 <= x_n_r_28; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_0_1 <= stage2_regs_r_9_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_0_2 <= stage2_regs_r_9_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_0_3 <= stage2_regs_r_9_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_0_4 <= stage2_regs_r_9_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_0_5 <= stage2_regs_r_9_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_0_6 <= stage2_regs_r_9_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_0_7 <= stage2_regs_r_9_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_0_8 <= stage2_regs_r_9_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_0_9 <= stage2_regs_r_9_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_0_10 <= stage2_regs_r_9_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_0_11 <= stage2_regs_r_9_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_9_1_0 <= a_2_r_28; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_1_1 <= stage2_regs_r_9_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_1_2 <= stage2_regs_r_9_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_1_3 <= stage2_regs_r_9_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_1_4 <= stage2_regs_r_9_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_1_5 <= stage2_regs_r_9_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_1_6 <= stage2_regs_r_9_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_1_7 <= stage2_regs_r_9_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_1_8 <= stage2_regs_r_9_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_1_9 <= stage2_regs_r_9_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_1_10 <= stage2_regs_r_9_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_9_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_9_1_11 <= stage2_regs_r_9_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_10_0_0 <= x_n_r_31; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_0_1 <= stage2_regs_r_10_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_0_2 <= stage2_regs_r_10_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_0_3 <= stage2_regs_r_10_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_0_4 <= stage2_regs_r_10_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_0_5 <= stage2_regs_r_10_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_0_6 <= stage2_regs_r_10_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_0_7 <= stage2_regs_r_10_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_0_8 <= stage2_regs_r_10_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_0_9 <= stage2_regs_r_10_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_0_10 <= stage2_regs_r_10_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_0_11 <= stage2_regs_r_10_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_10_1_0 <= a_2_r_31; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_1_1 <= stage2_regs_r_10_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_1_2 <= stage2_regs_r_10_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_1_3 <= stage2_regs_r_10_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_1_4 <= stage2_regs_r_10_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_1_5 <= stage2_regs_r_10_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_1_6 <= stage2_regs_r_10_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_1_7 <= stage2_regs_r_10_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_1_8 <= stage2_regs_r_10_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_1_9 <= stage2_regs_r_10_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_1_10 <= stage2_regs_r_10_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_10_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_10_1_11 <= stage2_regs_r_10_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_11_0_0 <= x_n_r_34; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_0_1 <= stage2_regs_r_11_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_0_2 <= stage2_regs_r_11_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_0_3 <= stage2_regs_r_11_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_0_4 <= stage2_regs_r_11_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_0_5 <= stage2_regs_r_11_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_0_6 <= stage2_regs_r_11_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_0_7 <= stage2_regs_r_11_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_0_8 <= stage2_regs_r_11_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_0_9 <= stage2_regs_r_11_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_0_10 <= stage2_regs_r_11_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_0_11 <= stage2_regs_r_11_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_11_1_0 <= a_2_r_34; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_1_1 <= stage2_regs_r_11_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_1_2 <= stage2_regs_r_11_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_1_3 <= stage2_regs_r_11_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_1_4 <= stage2_regs_r_11_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_1_5 <= stage2_regs_r_11_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_1_6 <= stage2_regs_r_11_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_1_7 <= stage2_regs_r_11_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_1_8 <= stage2_regs_r_11_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_1_9 <= stage2_regs_r_11_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_1_10 <= stage2_regs_r_11_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_11_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_11_1_11 <= stage2_regs_r_11_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_12_0_0 <= x_n_r_37; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_0_1 <= stage2_regs_r_12_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_0_2 <= stage2_regs_r_12_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_0_3 <= stage2_regs_r_12_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_0_4 <= stage2_regs_r_12_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_0_5 <= stage2_regs_r_12_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_0_6 <= stage2_regs_r_12_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_0_7 <= stage2_regs_r_12_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_0_8 <= stage2_regs_r_12_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_0_9 <= stage2_regs_r_12_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_0_10 <= stage2_regs_r_12_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_0_11 <= stage2_regs_r_12_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_12_1_0 <= a_2_r_37; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_1_1 <= stage2_regs_r_12_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_1_2 <= stage2_regs_r_12_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_1_3 <= stage2_regs_r_12_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_1_4 <= stage2_regs_r_12_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_1_5 <= stage2_regs_r_12_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_1_6 <= stage2_regs_r_12_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_1_7 <= stage2_regs_r_12_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_1_8 <= stage2_regs_r_12_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_1_9 <= stage2_regs_r_12_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_1_10 <= stage2_regs_r_12_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_12_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_12_1_11 <= stage2_regs_r_12_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_13_0_0 <= x_n_r_40; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_0_1 <= stage2_regs_r_13_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_0_2 <= stage2_regs_r_13_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_0_3 <= stage2_regs_r_13_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_0_4 <= stage2_regs_r_13_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_0_5 <= stage2_regs_r_13_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_0_6 <= stage2_regs_r_13_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_0_7 <= stage2_regs_r_13_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_0_8 <= stage2_regs_r_13_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_0_9 <= stage2_regs_r_13_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_0_10 <= stage2_regs_r_13_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_0_11 <= stage2_regs_r_13_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_13_1_0 <= a_2_r_40; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_1_1 <= stage2_regs_r_13_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_1_2 <= stage2_regs_r_13_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_1_3 <= stage2_regs_r_13_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_1_4 <= stage2_regs_r_13_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_1_5 <= stage2_regs_r_13_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_1_6 <= stage2_regs_r_13_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_1_7 <= stage2_regs_r_13_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_1_8 <= stage2_regs_r_13_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_1_9 <= stage2_regs_r_13_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_1_10 <= stage2_regs_r_13_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_13_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_13_1_11 <= stage2_regs_r_13_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_14_0_0 <= x_n_r_43; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_0_1 <= stage2_regs_r_14_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_0_2 <= stage2_regs_r_14_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_0_3 <= stage2_regs_r_14_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_0_4 <= stage2_regs_r_14_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_0_5 <= stage2_regs_r_14_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_0_6 <= stage2_regs_r_14_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_0_7 <= stage2_regs_r_14_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_0_8 <= stage2_regs_r_14_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_0_9 <= stage2_regs_r_14_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_0_10 <= stage2_regs_r_14_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_0_11 <= stage2_regs_r_14_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_14_1_0 <= a_2_r_43; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_1_1 <= stage2_regs_r_14_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_1_2 <= stage2_regs_r_14_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_1_3 <= stage2_regs_r_14_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_1_4 <= stage2_regs_r_14_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_1_5 <= stage2_regs_r_14_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_1_6 <= stage2_regs_r_14_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_1_7 <= stage2_regs_r_14_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_1_8 <= stage2_regs_r_14_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_1_9 <= stage2_regs_r_14_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_1_10 <= stage2_regs_r_14_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_14_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_14_1_11 <= stage2_regs_r_14_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_15_0_0 <= x_n_r_46; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_0_1 <= stage2_regs_r_15_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_0_2 <= stage2_regs_r_15_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_0_3 <= stage2_regs_r_15_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_0_4 <= stage2_regs_r_15_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_0_5 <= stage2_regs_r_15_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_0_6 <= stage2_regs_r_15_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_0_7 <= stage2_regs_r_15_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_0_8 <= stage2_regs_r_15_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_0_9 <= stage2_regs_r_15_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_0_10 <= stage2_regs_r_15_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_0_11 <= stage2_regs_r_15_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_15_1_0 <= a_2_r_46; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_1_1 <= stage2_regs_r_15_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_1_2 <= stage2_regs_r_15_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_1_3 <= stage2_regs_r_15_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_1_4 <= stage2_regs_r_15_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_1_5 <= stage2_regs_r_15_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_1_6 <= stage2_regs_r_15_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_1_7 <= stage2_regs_r_15_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_1_8 <= stage2_regs_r_15_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_1_9 <= stage2_regs_r_15_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_1_10 <= stage2_regs_r_15_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_15_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_15_1_11 <= stage2_regs_r_15_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_16_0_0 <= x_n_r_49; // @[FloatingPointDesigns.scala 2250:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_0_1 <= stage2_regs_r_16_0_0; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_0_2 <= stage2_regs_r_16_0_1; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_0_3 <= stage2_regs_r_16_0_2; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_0_4 <= stage2_regs_r_16_0_3; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_0_5 <= stage2_regs_r_16_0_4; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_0_6 <= stage2_regs_r_16_0_5; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_0_7 <= stage2_regs_r_16_0_6; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_0_8 <= stage2_regs_r_16_0_7; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_0_9 <= stage2_regs_r_16_0_8; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_0_10 <= stage2_regs_r_16_0_9; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_0_11 <= stage2_regs_r_16_0_10; // @[FloatingPointDesigns.scala 2214:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2247:26]
      stage2_regs_r_16_1_0 <= a_2_r_49; // @[FloatingPointDesigns.scala 2251:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_1_1 <= stage2_regs_r_16_1_0; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_1_2 <= stage2_regs_r_16_1_1; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_1_3 <= stage2_regs_r_16_1_2; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_1_4 <= stage2_regs_r_16_1_3; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_1_5 <= stage2_regs_r_16_1_4; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_1_6 <= stage2_regs_r_16_1_5; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_1_7 <= stage2_regs_r_16_1_6; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_1_8 <= stage2_regs_r_16_1_7; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_1_9 <= stage2_regs_r_16_1_8; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_1_10 <= stage2_regs_r_16_1_9; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2204:32]
      stage2_regs_r_16_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2204:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage2_regs_r_16_1_11 <= stage2_regs_r_16_1_10; // @[FloatingPointDesigns.scala 2215:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_0_1_0 <= a_2_r_2; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_0_1_1 <= stage3_regs_r_0_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_0_1_2 <= stage3_regs_r_0_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_0_1_3 <= stage3_regs_r_0_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_0_1_4 <= stage3_regs_r_0_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_0_1_5 <= stage3_regs_r_0_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_0_1_6 <= stage3_regs_r_0_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_0_1_7 <= stage3_regs_r_0_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_0_1_8 <= stage3_regs_r_0_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_1_1_0 <= a_2_r_5; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_1_1_1 <= stage3_regs_r_1_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_1_1_2 <= stage3_regs_r_1_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_1_1_3 <= stage3_regs_r_1_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_1_1_4 <= stage3_regs_r_1_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_1_1_5 <= stage3_regs_r_1_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_1_1_6 <= stage3_regs_r_1_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_1_1_7 <= stage3_regs_r_1_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_1_1_8 <= stage3_regs_r_1_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_2_1_0 <= a_2_r_8; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_2_1_1 <= stage3_regs_r_2_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_2_1_2 <= stage3_regs_r_2_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_2_1_3 <= stage3_regs_r_2_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_2_1_4 <= stage3_regs_r_2_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_2_1_5 <= stage3_regs_r_2_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_2_1_6 <= stage3_regs_r_2_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_2_1_7 <= stage3_regs_r_2_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_2_1_8 <= stage3_regs_r_2_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_3_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_3_1_0 <= a_2_r_11; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_3_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_3_1_1 <= stage3_regs_r_3_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_3_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_3_1_2 <= stage3_regs_r_3_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_3_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_3_1_3 <= stage3_regs_r_3_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_3_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_3_1_4 <= stage3_regs_r_3_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_3_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_3_1_5 <= stage3_regs_r_3_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_3_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_3_1_6 <= stage3_regs_r_3_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_3_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_3_1_7 <= stage3_regs_r_3_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_3_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_3_1_8 <= stage3_regs_r_3_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_4_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_4_1_0 <= a_2_r_14; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_4_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_4_1_1 <= stage3_regs_r_4_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_4_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_4_1_2 <= stage3_regs_r_4_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_4_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_4_1_3 <= stage3_regs_r_4_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_4_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_4_1_4 <= stage3_regs_r_4_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_4_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_4_1_5 <= stage3_regs_r_4_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_4_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_4_1_6 <= stage3_regs_r_4_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_4_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_4_1_7 <= stage3_regs_r_4_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_4_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_4_1_8 <= stage3_regs_r_4_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_5_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_5_1_0 <= a_2_r_17; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_5_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_5_1_1 <= stage3_regs_r_5_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_5_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_5_1_2 <= stage3_regs_r_5_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_5_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_5_1_3 <= stage3_regs_r_5_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_5_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_5_1_4 <= stage3_regs_r_5_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_5_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_5_1_5 <= stage3_regs_r_5_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_5_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_5_1_6 <= stage3_regs_r_5_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_5_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_5_1_7 <= stage3_regs_r_5_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_5_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_5_1_8 <= stage3_regs_r_5_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_6_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_6_1_0 <= a_2_r_20; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_6_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_6_1_1 <= stage3_regs_r_6_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_6_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_6_1_2 <= stage3_regs_r_6_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_6_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_6_1_3 <= stage3_regs_r_6_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_6_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_6_1_4 <= stage3_regs_r_6_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_6_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_6_1_5 <= stage3_regs_r_6_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_6_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_6_1_6 <= stage3_regs_r_6_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_6_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_6_1_7 <= stage3_regs_r_6_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_6_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_6_1_8 <= stage3_regs_r_6_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_7_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_7_1_0 <= a_2_r_23; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_7_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_7_1_1 <= stage3_regs_r_7_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_7_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_7_1_2 <= stage3_regs_r_7_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_7_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_7_1_3 <= stage3_regs_r_7_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_7_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_7_1_4 <= stage3_regs_r_7_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_7_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_7_1_5 <= stage3_regs_r_7_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_7_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_7_1_6 <= stage3_regs_r_7_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_7_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_7_1_7 <= stage3_regs_r_7_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_7_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_7_1_8 <= stage3_regs_r_7_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_8_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_8_1_0 <= a_2_r_26; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_8_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_8_1_1 <= stage3_regs_r_8_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_8_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_8_1_2 <= stage3_regs_r_8_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_8_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_8_1_3 <= stage3_regs_r_8_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_8_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_8_1_4 <= stage3_regs_r_8_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_8_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_8_1_5 <= stage3_regs_r_8_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_8_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_8_1_6 <= stage3_regs_r_8_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_8_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_8_1_7 <= stage3_regs_r_8_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_8_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_8_1_8 <= stage3_regs_r_8_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_9_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_9_1_0 <= a_2_r_29; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_9_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_9_1_1 <= stage3_regs_r_9_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_9_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_9_1_2 <= stage3_regs_r_9_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_9_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_9_1_3 <= stage3_regs_r_9_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_9_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_9_1_4 <= stage3_regs_r_9_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_9_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_9_1_5 <= stage3_regs_r_9_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_9_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_9_1_6 <= stage3_regs_r_9_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_9_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_9_1_7 <= stage3_regs_r_9_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_9_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_9_1_8 <= stage3_regs_r_9_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_10_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_10_1_0 <= a_2_r_32; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_10_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_10_1_1 <= stage3_regs_r_10_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_10_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_10_1_2 <= stage3_regs_r_10_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_10_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_10_1_3 <= stage3_regs_r_10_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_10_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_10_1_4 <= stage3_regs_r_10_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_10_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_10_1_5 <= stage3_regs_r_10_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_10_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_10_1_6 <= stage3_regs_r_10_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_10_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_10_1_7 <= stage3_regs_r_10_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_10_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_10_1_8 <= stage3_regs_r_10_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_11_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_11_1_0 <= a_2_r_35; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_11_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_11_1_1 <= stage3_regs_r_11_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_11_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_11_1_2 <= stage3_regs_r_11_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_11_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_11_1_3 <= stage3_regs_r_11_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_11_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_11_1_4 <= stage3_regs_r_11_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_11_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_11_1_5 <= stage3_regs_r_11_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_11_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_11_1_6 <= stage3_regs_r_11_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_11_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_11_1_7 <= stage3_regs_r_11_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_11_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_11_1_8 <= stage3_regs_r_11_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_12_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_12_1_0 <= a_2_r_38; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_12_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_12_1_1 <= stage3_regs_r_12_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_12_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_12_1_2 <= stage3_regs_r_12_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_12_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_12_1_3 <= stage3_regs_r_12_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_12_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_12_1_4 <= stage3_regs_r_12_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_12_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_12_1_5 <= stage3_regs_r_12_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_12_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_12_1_6 <= stage3_regs_r_12_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_12_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_12_1_7 <= stage3_regs_r_12_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_12_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_12_1_8 <= stage3_regs_r_12_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_13_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_13_1_0 <= a_2_r_41; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_13_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_13_1_1 <= stage3_regs_r_13_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_13_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_13_1_2 <= stage3_regs_r_13_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_13_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_13_1_3 <= stage3_regs_r_13_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_13_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_13_1_4 <= stage3_regs_r_13_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_13_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_13_1_5 <= stage3_regs_r_13_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_13_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_13_1_6 <= stage3_regs_r_13_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_13_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_13_1_7 <= stage3_regs_r_13_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_13_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_13_1_8 <= stage3_regs_r_13_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_14_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_14_1_0 <= a_2_r_44; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_14_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_14_1_1 <= stage3_regs_r_14_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_14_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_14_1_2 <= stage3_regs_r_14_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_14_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_14_1_3 <= stage3_regs_r_14_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_14_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_14_1_4 <= stage3_regs_r_14_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_14_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_14_1_5 <= stage3_regs_r_14_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_14_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_14_1_6 <= stage3_regs_r_14_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_14_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_14_1_7 <= stage3_regs_r_14_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_14_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_14_1_8 <= stage3_regs_r_14_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_15_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_15_1_0 <= a_2_r_47; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_15_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_15_1_1 <= stage3_regs_r_15_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_15_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_15_1_2 <= stage3_regs_r_15_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_15_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_15_1_3 <= stage3_regs_r_15_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_15_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_15_1_4 <= stage3_regs_r_15_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_15_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_15_1_5 <= stage3_regs_r_15_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_15_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_15_1_6 <= stage3_regs_r_15_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_15_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_15_1_7 <= stage3_regs_r_15_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_15_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_15_1_8 <= stage3_regs_r_15_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_16_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2256:26]
      stage3_regs_r_16_1_0 <= a_2_r_50; // @[FloatingPointDesigns.scala 2258:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_16_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_16_1_1 <= stage3_regs_r_16_1_0; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_16_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_16_1_2 <= stage3_regs_r_16_1_1; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_16_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_16_1_3 <= stage3_regs_r_16_1_2; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_16_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_16_1_4 <= stage3_regs_r_16_1_3; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_16_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_16_1_5 <= stage3_regs_r_16_1_4; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_16_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_16_1_6 <= stage3_regs_r_16_1_5; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_16_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_16_1_7 <= stage3_regs_r_16_1_6; // @[FloatingPointDesigns.scala 2219:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2205:32]
      stage3_regs_r_16_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2205:32]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2212:22]
      stage3_regs_r_16_1_8 <= stage3_regs_r_16_1_7; // @[FloatingPointDesigns.scala 2219:36]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  x_n_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  x_n_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  x_n_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  x_n_4 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  x_n_5 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  x_n_6 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  x_n_8 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  x_n_9 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  x_n_10 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  x_n_12 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  x_n_13 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  x_n_14 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  x_n_16 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  x_n_17 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  x_n_18 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  x_n_20 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  x_n_21 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  x_n_22 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  x_n_24 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  x_n_25 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  x_n_26 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  x_n_28 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  x_n_29 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  x_n_30 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  x_n_32 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  x_n_33 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  x_n_34 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  x_n_36 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  x_n_37 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  x_n_38 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  x_n_40 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  x_n_41 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  x_n_42 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  x_n_44 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  x_n_45 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  x_n_46 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  x_n_48 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  x_n_49 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  x_n_50 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  x_n_52 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  x_n_53 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  x_n_54 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  x_n_56 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  x_n_57 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  x_n_58 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  x_n_60 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  x_n_61 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  x_n_62 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  a_2_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  a_2_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  a_2_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  a_2_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  a_2_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  a_2_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  a_2_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  a_2_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  a_2_8 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  a_2_9 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  a_2_10 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  a_2_11 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  a_2_12 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  a_2_13 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  a_2_14 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  a_2_15 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  a_2_16 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  a_2_17 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  a_2_18 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  a_2_19 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  a_2_20 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  a_2_21 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  a_2_22 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  a_2_23 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  a_2_24 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  a_2_25 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  a_2_26 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  a_2_27 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  a_2_28 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  a_2_29 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  a_2_30 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  a_2_31 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  a_2_32 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  a_2_33 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  a_2_34 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  a_2_35 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  a_2_36 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  a_2_37 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  a_2_38 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  a_2_39 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  a_2_40 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  a_2_41 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  a_2_42 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  a_2_43 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  a_2_44 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  a_2_45 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  a_2_46 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  a_2_47 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  a_2_48 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  a_2_49 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  a_2_50 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  a_2_51 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  a_2_52 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  a_2_53 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  a_2_54 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  a_2_55 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  a_2_56 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  a_2_57 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  a_2_58 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  a_2_59 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  a_2_60 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  a_2_61 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  a_2_62 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  a_2_63 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  stage1_regs_0_0_0 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  stage1_regs_0_0_1 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  stage1_regs_0_0_2 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  stage1_regs_0_0_3 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  stage1_regs_0_0_4 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  stage1_regs_0_0_5 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  stage1_regs_0_0_6 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  stage1_regs_0_0_7 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  stage1_regs_0_0_8 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  stage1_regs_0_1_0 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  stage1_regs_0_1_1 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  stage1_regs_0_1_2 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  stage1_regs_0_1_3 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  stage1_regs_0_1_4 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  stage1_regs_0_1_5 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  stage1_regs_0_1_6 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  stage1_regs_0_1_7 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  stage1_regs_0_1_8 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  stage1_regs_1_0_0 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  stage1_regs_1_0_1 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  stage1_regs_1_0_2 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  stage1_regs_1_0_3 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  stage1_regs_1_0_4 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  stage1_regs_1_0_5 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  stage1_regs_1_0_6 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  stage1_regs_1_0_7 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  stage1_regs_1_0_8 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  stage1_regs_1_1_0 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  stage1_regs_1_1_1 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  stage1_regs_1_1_2 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  stage1_regs_1_1_3 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  stage1_regs_1_1_4 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  stage1_regs_1_1_5 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  stage1_regs_1_1_6 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  stage1_regs_1_1_7 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  stage1_regs_1_1_8 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  stage1_regs_2_0_0 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  stage1_regs_2_0_1 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  stage1_regs_2_0_2 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  stage1_regs_2_0_3 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  stage1_regs_2_0_4 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  stage1_regs_2_0_5 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  stage1_regs_2_0_6 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  stage1_regs_2_0_7 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  stage1_regs_2_0_8 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  stage1_regs_2_1_0 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  stage1_regs_2_1_1 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  stage1_regs_2_1_2 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  stage1_regs_2_1_3 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  stage1_regs_2_1_4 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  stage1_regs_2_1_5 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  stage1_regs_2_1_6 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  stage1_regs_2_1_7 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  stage1_regs_2_1_8 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  stage1_regs_3_0_0 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  stage1_regs_3_0_1 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  stage1_regs_3_0_2 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  stage1_regs_3_0_3 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  stage1_regs_3_0_4 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  stage1_regs_3_0_5 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  stage1_regs_3_0_6 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  stage1_regs_3_0_7 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  stage1_regs_3_0_8 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  stage1_regs_3_1_0 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  stage1_regs_3_1_1 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  stage1_regs_3_1_2 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  stage1_regs_3_1_3 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  stage1_regs_3_1_4 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  stage1_regs_3_1_5 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  stage1_regs_3_1_6 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  stage1_regs_3_1_7 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  stage1_regs_3_1_8 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  stage1_regs_4_0_0 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  stage1_regs_4_0_1 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  stage1_regs_4_0_2 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  stage1_regs_4_0_3 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  stage1_regs_4_0_4 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  stage1_regs_4_0_5 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  stage1_regs_4_0_6 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  stage1_regs_4_0_7 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  stage1_regs_4_0_8 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  stage1_regs_4_1_0 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  stage1_regs_4_1_1 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  stage1_regs_4_1_2 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  stage1_regs_4_1_3 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  stage1_regs_4_1_4 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  stage1_regs_4_1_5 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  stage1_regs_4_1_6 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  stage1_regs_4_1_7 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  stage1_regs_4_1_8 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  stage1_regs_5_0_0 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  stage1_regs_5_0_1 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  stage1_regs_5_0_2 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  stage1_regs_5_0_3 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  stage1_regs_5_0_4 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  stage1_regs_5_0_5 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  stage1_regs_5_0_6 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  stage1_regs_5_0_7 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  stage1_regs_5_0_8 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  stage1_regs_5_1_0 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  stage1_regs_5_1_1 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  stage1_regs_5_1_2 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  stage1_regs_5_1_3 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  stage1_regs_5_1_4 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  stage1_regs_5_1_5 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  stage1_regs_5_1_6 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  stage1_regs_5_1_7 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  stage1_regs_5_1_8 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  stage1_regs_6_0_0 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  stage1_regs_6_0_1 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  stage1_regs_6_0_2 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  stage1_regs_6_0_3 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  stage1_regs_6_0_4 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  stage1_regs_6_0_5 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  stage1_regs_6_0_6 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  stage1_regs_6_0_7 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  stage1_regs_6_0_8 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  stage1_regs_6_1_0 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  stage1_regs_6_1_1 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  stage1_regs_6_1_2 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  stage1_regs_6_1_3 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  stage1_regs_6_1_4 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  stage1_regs_6_1_5 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  stage1_regs_6_1_6 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  stage1_regs_6_1_7 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  stage1_regs_6_1_8 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  stage1_regs_7_0_0 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  stage1_regs_7_0_1 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  stage1_regs_7_0_2 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  stage1_regs_7_0_3 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  stage1_regs_7_0_4 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  stage1_regs_7_0_5 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  stage1_regs_7_0_6 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  stage1_regs_7_0_7 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  stage1_regs_7_0_8 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  stage1_regs_7_1_0 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  stage1_regs_7_1_1 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  stage1_regs_7_1_2 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  stage1_regs_7_1_3 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  stage1_regs_7_1_4 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  stage1_regs_7_1_5 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  stage1_regs_7_1_6 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  stage1_regs_7_1_7 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  stage1_regs_7_1_8 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  stage1_regs_8_0_0 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  stage1_regs_8_0_1 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  stage1_regs_8_0_2 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  stage1_regs_8_0_3 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  stage1_regs_8_0_4 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  stage1_regs_8_0_5 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  stage1_regs_8_0_6 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  stage1_regs_8_0_7 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  stage1_regs_8_0_8 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  stage1_regs_8_1_0 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  stage1_regs_8_1_1 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  stage1_regs_8_1_2 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  stage1_regs_8_1_3 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  stage1_regs_8_1_4 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  stage1_regs_8_1_5 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  stage1_regs_8_1_6 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  stage1_regs_8_1_7 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  stage1_regs_8_1_8 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  stage1_regs_9_0_0 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  stage1_regs_9_0_1 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  stage1_regs_9_0_2 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  stage1_regs_9_0_3 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  stage1_regs_9_0_4 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  stage1_regs_9_0_5 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  stage1_regs_9_0_6 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  stage1_regs_9_0_7 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  stage1_regs_9_0_8 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  stage1_regs_9_1_0 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  stage1_regs_9_1_1 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  stage1_regs_9_1_2 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  stage1_regs_9_1_3 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  stage1_regs_9_1_4 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  stage1_regs_9_1_5 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  stage1_regs_9_1_6 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  stage1_regs_9_1_7 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  stage1_regs_9_1_8 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  stage1_regs_10_0_0 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  stage1_regs_10_0_1 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  stage1_regs_10_0_2 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  stage1_regs_10_0_3 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  stage1_regs_10_0_4 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  stage1_regs_10_0_5 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  stage1_regs_10_0_6 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  stage1_regs_10_0_7 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  stage1_regs_10_0_8 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  stage1_regs_10_1_0 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  stage1_regs_10_1_1 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  stage1_regs_10_1_2 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  stage1_regs_10_1_3 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  stage1_regs_10_1_4 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  stage1_regs_10_1_5 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  stage1_regs_10_1_6 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  stage1_regs_10_1_7 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  stage1_regs_10_1_8 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  stage1_regs_11_0_0 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  stage1_regs_11_0_1 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  stage1_regs_11_0_2 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  stage1_regs_11_0_3 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  stage1_regs_11_0_4 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  stage1_regs_11_0_5 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  stage1_regs_11_0_6 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  stage1_regs_11_0_7 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  stage1_regs_11_0_8 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  stage1_regs_11_1_0 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  stage1_regs_11_1_1 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  stage1_regs_11_1_2 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  stage1_regs_11_1_3 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  stage1_regs_11_1_4 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  stage1_regs_11_1_5 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  stage1_regs_11_1_6 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  stage1_regs_11_1_7 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  stage1_regs_11_1_8 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  stage1_regs_12_0_0 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  stage1_regs_12_0_1 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  stage1_regs_12_0_2 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  stage1_regs_12_0_3 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  stage1_regs_12_0_4 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  stage1_regs_12_0_5 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  stage1_regs_12_0_6 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  stage1_regs_12_0_7 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  stage1_regs_12_0_8 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  stage1_regs_12_1_0 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  stage1_regs_12_1_1 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  stage1_regs_12_1_2 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  stage1_regs_12_1_3 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  stage1_regs_12_1_4 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  stage1_regs_12_1_5 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  stage1_regs_12_1_6 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  stage1_regs_12_1_7 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  stage1_regs_12_1_8 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  stage1_regs_13_0_0 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  stage1_regs_13_0_1 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  stage1_regs_13_0_2 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  stage1_regs_13_0_3 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  stage1_regs_13_0_4 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  stage1_regs_13_0_5 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  stage1_regs_13_0_6 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  stage1_regs_13_0_7 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  stage1_regs_13_0_8 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  stage1_regs_13_1_0 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  stage1_regs_13_1_1 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  stage1_regs_13_1_2 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  stage1_regs_13_1_3 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  stage1_regs_13_1_4 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  stage1_regs_13_1_5 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  stage1_regs_13_1_6 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  stage1_regs_13_1_7 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  stage1_regs_13_1_8 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  stage1_regs_14_0_0 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  stage1_regs_14_0_1 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  stage1_regs_14_0_2 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  stage1_regs_14_0_3 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  stage1_regs_14_0_4 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  stage1_regs_14_0_5 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  stage1_regs_14_0_6 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  stage1_regs_14_0_7 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  stage1_regs_14_0_8 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  stage1_regs_14_1_0 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  stage1_regs_14_1_1 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  stage1_regs_14_1_2 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  stage1_regs_14_1_3 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  stage1_regs_14_1_4 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  stage1_regs_14_1_5 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  stage1_regs_14_1_6 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  stage1_regs_14_1_7 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  stage1_regs_14_1_8 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  stage1_regs_15_0_0 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  stage1_regs_15_0_1 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  stage1_regs_15_0_2 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  stage1_regs_15_0_3 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  stage1_regs_15_0_4 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  stage1_regs_15_0_5 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  stage1_regs_15_0_6 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  stage1_regs_15_0_7 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  stage1_regs_15_0_8 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  stage1_regs_15_1_0 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  stage1_regs_15_1_1 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  stage1_regs_15_1_2 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  stage1_regs_15_1_3 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  stage1_regs_15_1_4 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  stage1_regs_15_1_5 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  stage1_regs_15_1_6 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  stage1_regs_15_1_7 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  stage1_regs_15_1_8 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  stage2_regs_0_0_0 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  stage2_regs_0_0_1 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  stage2_regs_0_0_2 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  stage2_regs_0_0_3 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  stage2_regs_0_0_4 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  stage2_regs_0_0_5 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  stage2_regs_0_0_6 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  stage2_regs_0_0_7 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  stage2_regs_0_0_8 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  stage2_regs_0_1_0 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  stage2_regs_0_1_1 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  stage2_regs_0_1_2 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  stage2_regs_0_1_3 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  stage2_regs_0_1_4 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  stage2_regs_0_1_5 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  stage2_regs_0_1_6 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  stage2_regs_0_1_7 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  stage2_regs_0_1_8 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  stage2_regs_1_0_0 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  stage2_regs_1_0_1 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  stage2_regs_1_0_2 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  stage2_regs_1_0_3 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  stage2_regs_1_0_4 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  stage2_regs_1_0_5 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  stage2_regs_1_0_6 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  stage2_regs_1_0_7 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  stage2_regs_1_0_8 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  stage2_regs_1_1_0 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  stage2_regs_1_1_1 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  stage2_regs_1_1_2 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  stage2_regs_1_1_3 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  stage2_regs_1_1_4 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  stage2_regs_1_1_5 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  stage2_regs_1_1_6 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  stage2_regs_1_1_7 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  stage2_regs_1_1_8 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  stage2_regs_2_0_0 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  stage2_regs_2_0_1 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  stage2_regs_2_0_2 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  stage2_regs_2_0_3 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  stage2_regs_2_0_4 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  stage2_regs_2_0_5 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  stage2_regs_2_0_6 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  stage2_regs_2_0_7 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  stage2_regs_2_0_8 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  stage2_regs_2_1_0 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  stage2_regs_2_1_1 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  stage2_regs_2_1_2 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  stage2_regs_2_1_3 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  stage2_regs_2_1_4 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  stage2_regs_2_1_5 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  stage2_regs_2_1_6 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  stage2_regs_2_1_7 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  stage2_regs_2_1_8 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  stage2_regs_3_0_0 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  stage2_regs_3_0_1 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  stage2_regs_3_0_2 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  stage2_regs_3_0_3 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  stage2_regs_3_0_4 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  stage2_regs_3_0_5 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  stage2_regs_3_0_6 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  stage2_regs_3_0_7 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  stage2_regs_3_0_8 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  stage2_regs_3_1_0 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  stage2_regs_3_1_1 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  stage2_regs_3_1_2 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  stage2_regs_3_1_3 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  stage2_regs_3_1_4 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  stage2_regs_3_1_5 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  stage2_regs_3_1_6 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  stage2_regs_3_1_7 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  stage2_regs_3_1_8 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  stage2_regs_4_0_0 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  stage2_regs_4_0_1 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  stage2_regs_4_0_2 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  stage2_regs_4_0_3 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  stage2_regs_4_0_4 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  stage2_regs_4_0_5 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  stage2_regs_4_0_6 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  stage2_regs_4_0_7 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  stage2_regs_4_0_8 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  stage2_regs_4_1_0 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  stage2_regs_4_1_1 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  stage2_regs_4_1_2 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  stage2_regs_4_1_3 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  stage2_regs_4_1_4 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  stage2_regs_4_1_5 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  stage2_regs_4_1_6 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  stage2_regs_4_1_7 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  stage2_regs_4_1_8 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  stage2_regs_5_0_0 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  stage2_regs_5_0_1 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  stage2_regs_5_0_2 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  stage2_regs_5_0_3 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  stage2_regs_5_0_4 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  stage2_regs_5_0_5 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  stage2_regs_5_0_6 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  stage2_regs_5_0_7 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  stage2_regs_5_0_8 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  stage2_regs_5_1_0 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  stage2_regs_5_1_1 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  stage2_regs_5_1_2 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  stage2_regs_5_1_3 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  stage2_regs_5_1_4 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  stage2_regs_5_1_5 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  stage2_regs_5_1_6 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  stage2_regs_5_1_7 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  stage2_regs_5_1_8 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  stage2_regs_6_0_0 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  stage2_regs_6_0_1 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  stage2_regs_6_0_2 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  stage2_regs_6_0_3 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  stage2_regs_6_0_4 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  stage2_regs_6_0_5 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  stage2_regs_6_0_6 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  stage2_regs_6_0_7 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  stage2_regs_6_0_8 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  stage2_regs_6_1_0 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  stage2_regs_6_1_1 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  stage2_regs_6_1_2 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  stage2_regs_6_1_3 = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  stage2_regs_6_1_4 = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  stage2_regs_6_1_5 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  stage2_regs_6_1_6 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  stage2_regs_6_1_7 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  stage2_regs_6_1_8 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  stage2_regs_7_0_0 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  stage2_regs_7_0_1 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  stage2_regs_7_0_2 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  stage2_regs_7_0_3 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  stage2_regs_7_0_4 = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  stage2_regs_7_0_5 = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  stage2_regs_7_0_6 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  stage2_regs_7_0_7 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  stage2_regs_7_0_8 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  stage2_regs_7_1_0 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  stage2_regs_7_1_1 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  stage2_regs_7_1_2 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  stage2_regs_7_1_3 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  stage2_regs_7_1_4 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  stage2_regs_7_1_5 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  stage2_regs_7_1_6 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  stage2_regs_7_1_7 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  stage2_regs_7_1_8 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  stage2_regs_8_0_0 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  stage2_regs_8_0_1 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  stage2_regs_8_0_2 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  stage2_regs_8_0_3 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  stage2_regs_8_0_4 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  stage2_regs_8_0_5 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  stage2_regs_8_0_6 = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  stage2_regs_8_0_7 = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  stage2_regs_8_0_8 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  stage2_regs_8_1_0 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  stage2_regs_8_1_1 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  stage2_regs_8_1_2 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  stage2_regs_8_1_3 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  stage2_regs_8_1_4 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  stage2_regs_8_1_5 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  stage2_regs_8_1_6 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  stage2_regs_8_1_7 = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  stage2_regs_8_1_8 = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  stage2_regs_9_0_0 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  stage2_regs_9_0_1 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  stage2_regs_9_0_2 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  stage2_regs_9_0_3 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  stage2_regs_9_0_4 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  stage2_regs_9_0_5 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  stage2_regs_9_0_6 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  stage2_regs_9_0_7 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  stage2_regs_9_0_8 = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  stage2_regs_9_1_0 = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  stage2_regs_9_1_1 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  stage2_regs_9_1_2 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  stage2_regs_9_1_3 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  stage2_regs_9_1_4 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  stage2_regs_9_1_5 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  stage2_regs_9_1_6 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  stage2_regs_9_1_7 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  stage2_regs_9_1_8 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  stage2_regs_10_0_0 = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  stage2_regs_10_0_1 = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  stage2_regs_10_0_2 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  stage2_regs_10_0_3 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  stage2_regs_10_0_4 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  stage2_regs_10_0_5 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  stage2_regs_10_0_6 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  stage2_regs_10_0_7 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  stage2_regs_10_0_8 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  stage2_regs_10_1_0 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  stage2_regs_10_1_1 = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  stage2_regs_10_1_2 = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  stage2_regs_10_1_3 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  stage2_regs_10_1_4 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  stage2_regs_10_1_5 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  stage2_regs_10_1_6 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  stage2_regs_10_1_7 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  stage2_regs_10_1_8 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  stage2_regs_11_0_0 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  stage2_regs_11_0_1 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  stage2_regs_11_0_2 = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  stage2_regs_11_0_3 = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  stage2_regs_11_0_4 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  stage2_regs_11_0_5 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  stage2_regs_11_0_6 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  stage2_regs_11_0_7 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  stage2_regs_11_0_8 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  stage2_regs_11_1_0 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  stage2_regs_11_1_1 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  stage2_regs_11_1_2 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  stage2_regs_11_1_3 = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  stage2_regs_11_1_4 = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  stage2_regs_11_1_5 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  stage2_regs_11_1_6 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  stage2_regs_11_1_7 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  stage2_regs_11_1_8 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  stage2_regs_12_0_0 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  stage2_regs_12_0_1 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  stage2_regs_12_0_2 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  stage2_regs_12_0_3 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  stage2_regs_12_0_4 = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  stage2_regs_12_0_5 = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  stage2_regs_12_0_6 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  stage2_regs_12_0_7 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  stage2_regs_12_0_8 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  stage2_regs_12_1_0 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  stage2_regs_12_1_1 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  stage2_regs_12_1_2 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  stage2_regs_12_1_3 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  stage2_regs_12_1_4 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  stage2_regs_12_1_5 = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  stage2_regs_12_1_6 = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  stage2_regs_12_1_7 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  stage2_regs_12_1_8 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  stage2_regs_13_0_0 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  stage2_regs_13_0_1 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  stage2_regs_13_0_2 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  stage2_regs_13_0_3 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  stage2_regs_13_0_4 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  stage2_regs_13_0_5 = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  stage2_regs_13_0_6 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  stage2_regs_13_0_7 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  stage2_regs_13_0_8 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  stage2_regs_13_1_0 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  stage2_regs_13_1_1 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  stage2_regs_13_1_2 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  stage2_regs_13_1_3 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  stage2_regs_13_1_4 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  stage2_regs_13_1_5 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  stage2_regs_13_1_6 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  stage2_regs_13_1_7 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  stage2_regs_13_1_8 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  stage2_regs_14_0_0 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  stage2_regs_14_0_1 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  stage2_regs_14_0_2 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  stage2_regs_14_0_3 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  stage2_regs_14_0_4 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  stage2_regs_14_0_5 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  stage2_regs_14_0_6 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  stage2_regs_14_0_7 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  stage2_regs_14_0_8 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  stage2_regs_14_1_0 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  stage2_regs_14_1_1 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  stage2_regs_14_1_2 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  stage2_regs_14_1_3 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  stage2_regs_14_1_4 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  stage2_regs_14_1_5 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  stage2_regs_14_1_6 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  stage2_regs_14_1_7 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  stage2_regs_14_1_8 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  stage2_regs_15_0_0 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  stage2_regs_15_0_1 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  stage2_regs_15_0_2 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  stage2_regs_15_0_3 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  stage2_regs_15_0_4 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  stage2_regs_15_0_5 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  stage2_regs_15_0_6 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  stage2_regs_15_0_7 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  stage2_regs_15_0_8 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  stage2_regs_15_1_0 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  stage2_regs_15_1_1 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  stage2_regs_15_1_2 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  stage2_regs_15_1_3 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  stage2_regs_15_1_4 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  stage2_regs_15_1_5 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  stage2_regs_15_1_6 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  stage2_regs_15_1_7 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  stage2_regs_15_1_8 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  stage3_regs_0_0_0 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  stage3_regs_0_0_1 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  stage3_regs_0_0_2 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  stage3_regs_0_0_3 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  stage3_regs_0_0_4 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  stage3_regs_0_0_5 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  stage3_regs_0_0_6 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  stage3_regs_0_0_7 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  stage3_regs_0_0_8 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  stage3_regs_0_0_9 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  stage3_regs_0_0_10 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  stage3_regs_0_0_11 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  stage3_regs_0_1_0 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  stage3_regs_0_1_1 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  stage3_regs_0_1_2 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  stage3_regs_0_1_3 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  stage3_regs_0_1_4 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  stage3_regs_0_1_5 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  stage3_regs_0_1_6 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  stage3_regs_0_1_7 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  stage3_regs_0_1_8 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  stage3_regs_0_1_9 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  stage3_regs_0_1_10 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  stage3_regs_0_1_11 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  stage3_regs_1_0_0 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  stage3_regs_1_0_1 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  stage3_regs_1_0_2 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  stage3_regs_1_0_3 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  stage3_regs_1_0_4 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  stage3_regs_1_0_5 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  stage3_regs_1_0_6 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  stage3_regs_1_0_7 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  stage3_regs_1_0_8 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  stage3_regs_1_0_9 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  stage3_regs_1_0_10 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  stage3_regs_1_0_11 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  stage3_regs_1_1_0 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  stage3_regs_1_1_1 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  stage3_regs_1_1_2 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  stage3_regs_1_1_3 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  stage3_regs_1_1_4 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  stage3_regs_1_1_5 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  stage3_regs_1_1_6 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  stage3_regs_1_1_7 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  stage3_regs_1_1_8 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  stage3_regs_1_1_9 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  stage3_regs_1_1_10 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  stage3_regs_1_1_11 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  stage3_regs_2_0_0 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  stage3_regs_2_0_1 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  stage3_regs_2_0_2 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  stage3_regs_2_0_3 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  stage3_regs_2_0_4 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  stage3_regs_2_0_5 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  stage3_regs_2_0_6 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  stage3_regs_2_0_7 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  stage3_regs_2_0_8 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  stage3_regs_2_0_9 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  stage3_regs_2_0_10 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  stage3_regs_2_0_11 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  stage3_regs_2_1_0 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  stage3_regs_2_1_1 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  stage3_regs_2_1_2 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  stage3_regs_2_1_3 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  stage3_regs_2_1_4 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  stage3_regs_2_1_5 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  stage3_regs_2_1_6 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  stage3_regs_2_1_7 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  stage3_regs_2_1_8 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  stage3_regs_2_1_9 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  stage3_regs_2_1_10 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  stage3_regs_2_1_11 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  stage3_regs_3_0_0 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  stage3_regs_3_0_1 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  stage3_regs_3_0_2 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  stage3_regs_3_0_3 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  stage3_regs_3_0_4 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  stage3_regs_3_0_5 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  stage3_regs_3_0_6 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  stage3_regs_3_0_7 = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  stage3_regs_3_0_8 = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  stage3_regs_3_0_9 = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  stage3_regs_3_0_10 = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  stage3_regs_3_0_11 = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  stage3_regs_3_1_0 = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  stage3_regs_3_1_1 = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  stage3_regs_3_1_2 = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  stage3_regs_3_1_3 = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  stage3_regs_3_1_4 = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  stage3_regs_3_1_5 = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  stage3_regs_3_1_6 = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  stage3_regs_3_1_7 = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  stage3_regs_3_1_8 = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  stage3_regs_3_1_9 = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  stage3_regs_3_1_10 = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  stage3_regs_3_1_11 = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  stage3_regs_4_0_0 = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  stage3_regs_4_0_1 = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  stage3_regs_4_0_2 = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  stage3_regs_4_0_3 = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  stage3_regs_4_0_4 = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  stage3_regs_4_0_5 = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  stage3_regs_4_0_6 = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  stage3_regs_4_0_7 = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  stage3_regs_4_0_8 = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  stage3_regs_4_0_9 = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  stage3_regs_4_0_10 = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  stage3_regs_4_0_11 = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  stage3_regs_4_1_0 = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  stage3_regs_4_1_1 = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  stage3_regs_4_1_2 = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  stage3_regs_4_1_3 = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  stage3_regs_4_1_4 = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  stage3_regs_4_1_5 = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  stage3_regs_4_1_6 = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  stage3_regs_4_1_7 = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  stage3_regs_4_1_8 = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  stage3_regs_4_1_9 = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  stage3_regs_4_1_10 = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  stage3_regs_4_1_11 = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  stage3_regs_5_0_0 = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  stage3_regs_5_0_1 = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  stage3_regs_5_0_2 = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  stage3_regs_5_0_3 = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  stage3_regs_5_0_4 = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  stage3_regs_5_0_5 = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  stage3_regs_5_0_6 = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  stage3_regs_5_0_7 = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  stage3_regs_5_0_8 = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  stage3_regs_5_0_9 = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  stage3_regs_5_0_10 = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  stage3_regs_5_0_11 = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  stage3_regs_5_1_0 = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  stage3_regs_5_1_1 = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  stage3_regs_5_1_2 = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  stage3_regs_5_1_3 = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  stage3_regs_5_1_4 = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  stage3_regs_5_1_5 = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  stage3_regs_5_1_6 = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  stage3_regs_5_1_7 = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  stage3_regs_5_1_8 = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  stage3_regs_5_1_9 = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  stage3_regs_5_1_10 = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  stage3_regs_5_1_11 = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  stage3_regs_6_0_0 = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  stage3_regs_6_0_1 = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  stage3_regs_6_0_2 = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  stage3_regs_6_0_3 = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  stage3_regs_6_0_4 = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  stage3_regs_6_0_5 = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  stage3_regs_6_0_6 = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  stage3_regs_6_0_7 = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  stage3_regs_6_0_8 = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  stage3_regs_6_0_9 = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  stage3_regs_6_0_10 = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  stage3_regs_6_0_11 = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  stage3_regs_6_1_0 = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  stage3_regs_6_1_1 = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  stage3_regs_6_1_2 = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  stage3_regs_6_1_3 = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  stage3_regs_6_1_4 = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  stage3_regs_6_1_5 = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  stage3_regs_6_1_6 = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  stage3_regs_6_1_7 = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  stage3_regs_6_1_8 = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  stage3_regs_6_1_9 = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  stage3_regs_6_1_10 = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  stage3_regs_6_1_11 = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  stage3_regs_7_0_0 = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  stage3_regs_7_0_1 = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  stage3_regs_7_0_2 = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  stage3_regs_7_0_3 = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  stage3_regs_7_0_4 = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  stage3_regs_7_0_5 = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  stage3_regs_7_0_6 = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  stage3_regs_7_0_7 = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  stage3_regs_7_0_8 = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  stage3_regs_7_0_9 = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  stage3_regs_7_0_10 = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  stage3_regs_7_0_11 = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  stage3_regs_7_1_0 = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  stage3_regs_7_1_1 = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  stage3_regs_7_1_2 = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  stage3_regs_7_1_3 = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  stage3_regs_7_1_4 = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  stage3_regs_7_1_5 = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  stage3_regs_7_1_6 = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  stage3_regs_7_1_7 = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  stage3_regs_7_1_8 = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  stage3_regs_7_1_9 = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  stage3_regs_7_1_10 = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  stage3_regs_7_1_11 = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  stage3_regs_8_0_0 = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  stage3_regs_8_0_1 = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  stage3_regs_8_0_2 = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  stage3_regs_8_0_3 = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  stage3_regs_8_0_4 = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  stage3_regs_8_0_5 = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  stage3_regs_8_0_6 = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  stage3_regs_8_0_7 = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  stage3_regs_8_0_8 = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  stage3_regs_8_0_9 = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  stage3_regs_8_0_10 = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  stage3_regs_8_0_11 = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  stage3_regs_8_1_0 = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  stage3_regs_8_1_1 = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  stage3_regs_8_1_2 = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  stage3_regs_8_1_3 = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  stage3_regs_8_1_4 = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  stage3_regs_8_1_5 = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  stage3_regs_8_1_6 = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  stage3_regs_8_1_7 = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  stage3_regs_8_1_8 = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  stage3_regs_8_1_9 = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  stage3_regs_8_1_10 = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  stage3_regs_8_1_11 = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  stage3_regs_9_0_0 = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  stage3_regs_9_0_1 = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  stage3_regs_9_0_2 = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  stage3_regs_9_0_3 = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  stage3_regs_9_0_4 = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  stage3_regs_9_0_5 = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  stage3_regs_9_0_6 = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  stage3_regs_9_0_7 = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  stage3_regs_9_0_8 = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  stage3_regs_9_0_9 = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  stage3_regs_9_0_10 = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  stage3_regs_9_0_11 = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  stage3_regs_9_1_0 = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  stage3_regs_9_1_1 = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  stage3_regs_9_1_2 = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  stage3_regs_9_1_3 = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  stage3_regs_9_1_4 = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  stage3_regs_9_1_5 = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  stage3_regs_9_1_6 = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  stage3_regs_9_1_7 = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  stage3_regs_9_1_8 = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  stage3_regs_9_1_9 = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  stage3_regs_9_1_10 = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  stage3_regs_9_1_11 = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  stage3_regs_10_0_0 = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  stage3_regs_10_0_1 = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  stage3_regs_10_0_2 = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  stage3_regs_10_0_3 = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  stage3_regs_10_0_4 = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  stage3_regs_10_0_5 = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  stage3_regs_10_0_6 = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  stage3_regs_10_0_7 = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  stage3_regs_10_0_8 = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  stage3_regs_10_0_9 = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  stage3_regs_10_0_10 = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  stage3_regs_10_0_11 = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  stage3_regs_10_1_0 = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  stage3_regs_10_1_1 = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  stage3_regs_10_1_2 = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  stage3_regs_10_1_3 = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  stage3_regs_10_1_4 = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  stage3_regs_10_1_5 = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  stage3_regs_10_1_6 = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  stage3_regs_10_1_7 = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  stage3_regs_10_1_8 = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  stage3_regs_10_1_9 = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  stage3_regs_10_1_10 = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  stage3_regs_10_1_11 = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  stage3_regs_11_0_0 = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  stage3_regs_11_0_1 = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  stage3_regs_11_0_2 = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  stage3_regs_11_0_3 = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  stage3_regs_11_0_4 = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  stage3_regs_11_0_5 = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  stage3_regs_11_0_6 = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  stage3_regs_11_0_7 = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  stage3_regs_11_0_8 = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  stage3_regs_11_0_9 = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  stage3_regs_11_0_10 = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  stage3_regs_11_0_11 = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  stage3_regs_11_1_0 = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  stage3_regs_11_1_1 = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  stage3_regs_11_1_2 = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  stage3_regs_11_1_3 = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  stage3_regs_11_1_4 = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  stage3_regs_11_1_5 = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  stage3_regs_11_1_6 = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  stage3_regs_11_1_7 = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  stage3_regs_11_1_8 = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  stage3_regs_11_1_9 = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  stage3_regs_11_1_10 = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  stage3_regs_11_1_11 = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  stage3_regs_12_0_0 = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  stage3_regs_12_0_1 = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  stage3_regs_12_0_2 = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  stage3_regs_12_0_3 = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  stage3_regs_12_0_4 = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  stage3_regs_12_0_5 = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  stage3_regs_12_0_6 = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  stage3_regs_12_0_7 = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  stage3_regs_12_0_8 = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  stage3_regs_12_0_9 = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  stage3_regs_12_0_10 = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  stage3_regs_12_0_11 = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  stage3_regs_12_1_0 = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  stage3_regs_12_1_1 = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  stage3_regs_12_1_2 = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  stage3_regs_12_1_3 = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  stage3_regs_12_1_4 = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  stage3_regs_12_1_5 = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  stage3_regs_12_1_6 = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  stage3_regs_12_1_7 = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  stage3_regs_12_1_8 = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  stage3_regs_12_1_9 = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  stage3_regs_12_1_10 = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  stage3_regs_12_1_11 = _RAND_999[31:0];
  _RAND_1000 = {1{`RANDOM}};
  stage3_regs_13_0_0 = _RAND_1000[31:0];
  _RAND_1001 = {1{`RANDOM}};
  stage3_regs_13_0_1 = _RAND_1001[31:0];
  _RAND_1002 = {1{`RANDOM}};
  stage3_regs_13_0_2 = _RAND_1002[31:0];
  _RAND_1003 = {1{`RANDOM}};
  stage3_regs_13_0_3 = _RAND_1003[31:0];
  _RAND_1004 = {1{`RANDOM}};
  stage3_regs_13_0_4 = _RAND_1004[31:0];
  _RAND_1005 = {1{`RANDOM}};
  stage3_regs_13_0_5 = _RAND_1005[31:0];
  _RAND_1006 = {1{`RANDOM}};
  stage3_regs_13_0_6 = _RAND_1006[31:0];
  _RAND_1007 = {1{`RANDOM}};
  stage3_regs_13_0_7 = _RAND_1007[31:0];
  _RAND_1008 = {1{`RANDOM}};
  stage3_regs_13_0_8 = _RAND_1008[31:0];
  _RAND_1009 = {1{`RANDOM}};
  stage3_regs_13_0_9 = _RAND_1009[31:0];
  _RAND_1010 = {1{`RANDOM}};
  stage3_regs_13_0_10 = _RAND_1010[31:0];
  _RAND_1011 = {1{`RANDOM}};
  stage3_regs_13_0_11 = _RAND_1011[31:0];
  _RAND_1012 = {1{`RANDOM}};
  stage3_regs_13_1_0 = _RAND_1012[31:0];
  _RAND_1013 = {1{`RANDOM}};
  stage3_regs_13_1_1 = _RAND_1013[31:0];
  _RAND_1014 = {1{`RANDOM}};
  stage3_regs_13_1_2 = _RAND_1014[31:0];
  _RAND_1015 = {1{`RANDOM}};
  stage3_regs_13_1_3 = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  stage3_regs_13_1_4 = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  stage3_regs_13_1_5 = _RAND_1017[31:0];
  _RAND_1018 = {1{`RANDOM}};
  stage3_regs_13_1_6 = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  stage3_regs_13_1_7 = _RAND_1019[31:0];
  _RAND_1020 = {1{`RANDOM}};
  stage3_regs_13_1_8 = _RAND_1020[31:0];
  _RAND_1021 = {1{`RANDOM}};
  stage3_regs_13_1_9 = _RAND_1021[31:0];
  _RAND_1022 = {1{`RANDOM}};
  stage3_regs_13_1_10 = _RAND_1022[31:0];
  _RAND_1023 = {1{`RANDOM}};
  stage3_regs_13_1_11 = _RAND_1023[31:0];
  _RAND_1024 = {1{`RANDOM}};
  stage3_regs_14_0_0 = _RAND_1024[31:0];
  _RAND_1025 = {1{`RANDOM}};
  stage3_regs_14_0_1 = _RAND_1025[31:0];
  _RAND_1026 = {1{`RANDOM}};
  stage3_regs_14_0_2 = _RAND_1026[31:0];
  _RAND_1027 = {1{`RANDOM}};
  stage3_regs_14_0_3 = _RAND_1027[31:0];
  _RAND_1028 = {1{`RANDOM}};
  stage3_regs_14_0_4 = _RAND_1028[31:0];
  _RAND_1029 = {1{`RANDOM}};
  stage3_regs_14_0_5 = _RAND_1029[31:0];
  _RAND_1030 = {1{`RANDOM}};
  stage3_regs_14_0_6 = _RAND_1030[31:0];
  _RAND_1031 = {1{`RANDOM}};
  stage3_regs_14_0_7 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  stage3_regs_14_0_8 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  stage3_regs_14_0_9 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  stage3_regs_14_0_10 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  stage3_regs_14_0_11 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  stage3_regs_14_1_0 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  stage3_regs_14_1_1 = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  stage3_regs_14_1_2 = _RAND_1038[31:0];
  _RAND_1039 = {1{`RANDOM}};
  stage3_regs_14_1_3 = _RAND_1039[31:0];
  _RAND_1040 = {1{`RANDOM}};
  stage3_regs_14_1_4 = _RAND_1040[31:0];
  _RAND_1041 = {1{`RANDOM}};
  stage3_regs_14_1_5 = _RAND_1041[31:0];
  _RAND_1042 = {1{`RANDOM}};
  stage3_regs_14_1_6 = _RAND_1042[31:0];
  _RAND_1043 = {1{`RANDOM}};
  stage3_regs_14_1_7 = _RAND_1043[31:0];
  _RAND_1044 = {1{`RANDOM}};
  stage3_regs_14_1_8 = _RAND_1044[31:0];
  _RAND_1045 = {1{`RANDOM}};
  stage3_regs_14_1_9 = _RAND_1045[31:0];
  _RAND_1046 = {1{`RANDOM}};
  stage3_regs_14_1_10 = _RAND_1046[31:0];
  _RAND_1047 = {1{`RANDOM}};
  stage3_regs_14_1_11 = _RAND_1047[31:0];
  _RAND_1048 = {1{`RANDOM}};
  stage3_regs_15_0_0 = _RAND_1048[31:0];
  _RAND_1049 = {1{`RANDOM}};
  stage3_regs_15_0_1 = _RAND_1049[31:0];
  _RAND_1050 = {1{`RANDOM}};
  stage3_regs_15_0_2 = _RAND_1050[31:0];
  _RAND_1051 = {1{`RANDOM}};
  stage3_regs_15_0_3 = _RAND_1051[31:0];
  _RAND_1052 = {1{`RANDOM}};
  stage3_regs_15_0_4 = _RAND_1052[31:0];
  _RAND_1053 = {1{`RANDOM}};
  stage3_regs_15_0_5 = _RAND_1053[31:0];
  _RAND_1054 = {1{`RANDOM}};
  stage3_regs_15_0_6 = _RAND_1054[31:0];
  _RAND_1055 = {1{`RANDOM}};
  stage3_regs_15_0_7 = _RAND_1055[31:0];
  _RAND_1056 = {1{`RANDOM}};
  stage3_regs_15_0_8 = _RAND_1056[31:0];
  _RAND_1057 = {1{`RANDOM}};
  stage3_regs_15_0_9 = _RAND_1057[31:0];
  _RAND_1058 = {1{`RANDOM}};
  stage3_regs_15_0_10 = _RAND_1058[31:0];
  _RAND_1059 = {1{`RANDOM}};
  stage3_regs_15_0_11 = _RAND_1059[31:0];
  _RAND_1060 = {1{`RANDOM}};
  stage3_regs_15_1_0 = _RAND_1060[31:0];
  _RAND_1061 = {1{`RANDOM}};
  stage3_regs_15_1_1 = _RAND_1061[31:0];
  _RAND_1062 = {1{`RANDOM}};
  stage3_regs_15_1_2 = _RAND_1062[31:0];
  _RAND_1063 = {1{`RANDOM}};
  stage3_regs_15_1_3 = _RAND_1063[31:0];
  _RAND_1064 = {1{`RANDOM}};
  stage3_regs_15_1_4 = _RAND_1064[31:0];
  _RAND_1065 = {1{`RANDOM}};
  stage3_regs_15_1_5 = _RAND_1065[31:0];
  _RAND_1066 = {1{`RANDOM}};
  stage3_regs_15_1_6 = _RAND_1066[31:0];
  _RAND_1067 = {1{`RANDOM}};
  stage3_regs_15_1_7 = _RAND_1067[31:0];
  _RAND_1068 = {1{`RANDOM}};
  stage3_regs_15_1_8 = _RAND_1068[31:0];
  _RAND_1069 = {1{`RANDOM}};
  stage3_regs_15_1_9 = _RAND_1069[31:0];
  _RAND_1070 = {1{`RANDOM}};
  stage3_regs_15_1_10 = _RAND_1070[31:0];
  _RAND_1071 = {1{`RANDOM}};
  stage3_regs_15_1_11 = _RAND_1071[31:0];
  _RAND_1072 = {1{`RANDOM}};
  stage4_regs_0_1_0 = _RAND_1072[31:0];
  _RAND_1073 = {1{`RANDOM}};
  stage4_regs_0_1_1 = _RAND_1073[31:0];
  _RAND_1074 = {1{`RANDOM}};
  stage4_regs_0_1_2 = _RAND_1074[31:0];
  _RAND_1075 = {1{`RANDOM}};
  stage4_regs_0_1_3 = _RAND_1075[31:0];
  _RAND_1076 = {1{`RANDOM}};
  stage4_regs_0_1_4 = _RAND_1076[31:0];
  _RAND_1077 = {1{`RANDOM}};
  stage4_regs_0_1_5 = _RAND_1077[31:0];
  _RAND_1078 = {1{`RANDOM}};
  stage4_regs_0_1_6 = _RAND_1078[31:0];
  _RAND_1079 = {1{`RANDOM}};
  stage4_regs_0_1_7 = _RAND_1079[31:0];
  _RAND_1080 = {1{`RANDOM}};
  stage4_regs_0_1_8 = _RAND_1080[31:0];
  _RAND_1081 = {1{`RANDOM}};
  stage4_regs_1_1_0 = _RAND_1081[31:0];
  _RAND_1082 = {1{`RANDOM}};
  stage4_regs_1_1_1 = _RAND_1082[31:0];
  _RAND_1083 = {1{`RANDOM}};
  stage4_regs_1_1_2 = _RAND_1083[31:0];
  _RAND_1084 = {1{`RANDOM}};
  stage4_regs_1_1_3 = _RAND_1084[31:0];
  _RAND_1085 = {1{`RANDOM}};
  stage4_regs_1_1_4 = _RAND_1085[31:0];
  _RAND_1086 = {1{`RANDOM}};
  stage4_regs_1_1_5 = _RAND_1086[31:0];
  _RAND_1087 = {1{`RANDOM}};
  stage4_regs_1_1_6 = _RAND_1087[31:0];
  _RAND_1088 = {1{`RANDOM}};
  stage4_regs_1_1_7 = _RAND_1088[31:0];
  _RAND_1089 = {1{`RANDOM}};
  stage4_regs_1_1_8 = _RAND_1089[31:0];
  _RAND_1090 = {1{`RANDOM}};
  stage4_regs_2_1_0 = _RAND_1090[31:0];
  _RAND_1091 = {1{`RANDOM}};
  stage4_regs_2_1_1 = _RAND_1091[31:0];
  _RAND_1092 = {1{`RANDOM}};
  stage4_regs_2_1_2 = _RAND_1092[31:0];
  _RAND_1093 = {1{`RANDOM}};
  stage4_regs_2_1_3 = _RAND_1093[31:0];
  _RAND_1094 = {1{`RANDOM}};
  stage4_regs_2_1_4 = _RAND_1094[31:0];
  _RAND_1095 = {1{`RANDOM}};
  stage4_regs_2_1_5 = _RAND_1095[31:0];
  _RAND_1096 = {1{`RANDOM}};
  stage4_regs_2_1_6 = _RAND_1096[31:0];
  _RAND_1097 = {1{`RANDOM}};
  stage4_regs_2_1_7 = _RAND_1097[31:0];
  _RAND_1098 = {1{`RANDOM}};
  stage4_regs_2_1_8 = _RAND_1098[31:0];
  _RAND_1099 = {1{`RANDOM}};
  stage4_regs_3_1_0 = _RAND_1099[31:0];
  _RAND_1100 = {1{`RANDOM}};
  stage4_regs_3_1_1 = _RAND_1100[31:0];
  _RAND_1101 = {1{`RANDOM}};
  stage4_regs_3_1_2 = _RAND_1101[31:0];
  _RAND_1102 = {1{`RANDOM}};
  stage4_regs_3_1_3 = _RAND_1102[31:0];
  _RAND_1103 = {1{`RANDOM}};
  stage4_regs_3_1_4 = _RAND_1103[31:0];
  _RAND_1104 = {1{`RANDOM}};
  stage4_regs_3_1_5 = _RAND_1104[31:0];
  _RAND_1105 = {1{`RANDOM}};
  stage4_regs_3_1_6 = _RAND_1105[31:0];
  _RAND_1106 = {1{`RANDOM}};
  stage4_regs_3_1_7 = _RAND_1106[31:0];
  _RAND_1107 = {1{`RANDOM}};
  stage4_regs_3_1_8 = _RAND_1107[31:0];
  _RAND_1108 = {1{`RANDOM}};
  stage4_regs_4_1_0 = _RAND_1108[31:0];
  _RAND_1109 = {1{`RANDOM}};
  stage4_regs_4_1_1 = _RAND_1109[31:0];
  _RAND_1110 = {1{`RANDOM}};
  stage4_regs_4_1_2 = _RAND_1110[31:0];
  _RAND_1111 = {1{`RANDOM}};
  stage4_regs_4_1_3 = _RAND_1111[31:0];
  _RAND_1112 = {1{`RANDOM}};
  stage4_regs_4_1_4 = _RAND_1112[31:0];
  _RAND_1113 = {1{`RANDOM}};
  stage4_regs_4_1_5 = _RAND_1113[31:0];
  _RAND_1114 = {1{`RANDOM}};
  stage4_regs_4_1_6 = _RAND_1114[31:0];
  _RAND_1115 = {1{`RANDOM}};
  stage4_regs_4_1_7 = _RAND_1115[31:0];
  _RAND_1116 = {1{`RANDOM}};
  stage4_regs_4_1_8 = _RAND_1116[31:0];
  _RAND_1117 = {1{`RANDOM}};
  stage4_regs_5_1_0 = _RAND_1117[31:0];
  _RAND_1118 = {1{`RANDOM}};
  stage4_regs_5_1_1 = _RAND_1118[31:0];
  _RAND_1119 = {1{`RANDOM}};
  stage4_regs_5_1_2 = _RAND_1119[31:0];
  _RAND_1120 = {1{`RANDOM}};
  stage4_regs_5_1_3 = _RAND_1120[31:0];
  _RAND_1121 = {1{`RANDOM}};
  stage4_regs_5_1_4 = _RAND_1121[31:0];
  _RAND_1122 = {1{`RANDOM}};
  stage4_regs_5_1_5 = _RAND_1122[31:0];
  _RAND_1123 = {1{`RANDOM}};
  stage4_regs_5_1_6 = _RAND_1123[31:0];
  _RAND_1124 = {1{`RANDOM}};
  stage4_regs_5_1_7 = _RAND_1124[31:0];
  _RAND_1125 = {1{`RANDOM}};
  stage4_regs_5_1_8 = _RAND_1125[31:0];
  _RAND_1126 = {1{`RANDOM}};
  stage4_regs_6_1_0 = _RAND_1126[31:0];
  _RAND_1127 = {1{`RANDOM}};
  stage4_regs_6_1_1 = _RAND_1127[31:0];
  _RAND_1128 = {1{`RANDOM}};
  stage4_regs_6_1_2 = _RAND_1128[31:0];
  _RAND_1129 = {1{`RANDOM}};
  stage4_regs_6_1_3 = _RAND_1129[31:0];
  _RAND_1130 = {1{`RANDOM}};
  stage4_regs_6_1_4 = _RAND_1130[31:0];
  _RAND_1131 = {1{`RANDOM}};
  stage4_regs_6_1_5 = _RAND_1131[31:0];
  _RAND_1132 = {1{`RANDOM}};
  stage4_regs_6_1_6 = _RAND_1132[31:0];
  _RAND_1133 = {1{`RANDOM}};
  stage4_regs_6_1_7 = _RAND_1133[31:0];
  _RAND_1134 = {1{`RANDOM}};
  stage4_regs_6_1_8 = _RAND_1134[31:0];
  _RAND_1135 = {1{`RANDOM}};
  stage4_regs_7_1_0 = _RAND_1135[31:0];
  _RAND_1136 = {1{`RANDOM}};
  stage4_regs_7_1_1 = _RAND_1136[31:0];
  _RAND_1137 = {1{`RANDOM}};
  stage4_regs_7_1_2 = _RAND_1137[31:0];
  _RAND_1138 = {1{`RANDOM}};
  stage4_regs_7_1_3 = _RAND_1138[31:0];
  _RAND_1139 = {1{`RANDOM}};
  stage4_regs_7_1_4 = _RAND_1139[31:0];
  _RAND_1140 = {1{`RANDOM}};
  stage4_regs_7_1_5 = _RAND_1140[31:0];
  _RAND_1141 = {1{`RANDOM}};
  stage4_regs_7_1_6 = _RAND_1141[31:0];
  _RAND_1142 = {1{`RANDOM}};
  stage4_regs_7_1_7 = _RAND_1142[31:0];
  _RAND_1143 = {1{`RANDOM}};
  stage4_regs_7_1_8 = _RAND_1143[31:0];
  _RAND_1144 = {1{`RANDOM}};
  stage4_regs_8_1_0 = _RAND_1144[31:0];
  _RAND_1145 = {1{`RANDOM}};
  stage4_regs_8_1_1 = _RAND_1145[31:0];
  _RAND_1146 = {1{`RANDOM}};
  stage4_regs_8_1_2 = _RAND_1146[31:0];
  _RAND_1147 = {1{`RANDOM}};
  stage4_regs_8_1_3 = _RAND_1147[31:0];
  _RAND_1148 = {1{`RANDOM}};
  stage4_regs_8_1_4 = _RAND_1148[31:0];
  _RAND_1149 = {1{`RANDOM}};
  stage4_regs_8_1_5 = _RAND_1149[31:0];
  _RAND_1150 = {1{`RANDOM}};
  stage4_regs_8_1_6 = _RAND_1150[31:0];
  _RAND_1151 = {1{`RANDOM}};
  stage4_regs_8_1_7 = _RAND_1151[31:0];
  _RAND_1152 = {1{`RANDOM}};
  stage4_regs_8_1_8 = _RAND_1152[31:0];
  _RAND_1153 = {1{`RANDOM}};
  stage4_regs_9_1_0 = _RAND_1153[31:0];
  _RAND_1154 = {1{`RANDOM}};
  stage4_regs_9_1_1 = _RAND_1154[31:0];
  _RAND_1155 = {1{`RANDOM}};
  stage4_regs_9_1_2 = _RAND_1155[31:0];
  _RAND_1156 = {1{`RANDOM}};
  stage4_regs_9_1_3 = _RAND_1156[31:0];
  _RAND_1157 = {1{`RANDOM}};
  stage4_regs_9_1_4 = _RAND_1157[31:0];
  _RAND_1158 = {1{`RANDOM}};
  stage4_regs_9_1_5 = _RAND_1158[31:0];
  _RAND_1159 = {1{`RANDOM}};
  stage4_regs_9_1_6 = _RAND_1159[31:0];
  _RAND_1160 = {1{`RANDOM}};
  stage4_regs_9_1_7 = _RAND_1160[31:0];
  _RAND_1161 = {1{`RANDOM}};
  stage4_regs_9_1_8 = _RAND_1161[31:0];
  _RAND_1162 = {1{`RANDOM}};
  stage4_regs_10_1_0 = _RAND_1162[31:0];
  _RAND_1163 = {1{`RANDOM}};
  stage4_regs_10_1_1 = _RAND_1163[31:0];
  _RAND_1164 = {1{`RANDOM}};
  stage4_regs_10_1_2 = _RAND_1164[31:0];
  _RAND_1165 = {1{`RANDOM}};
  stage4_regs_10_1_3 = _RAND_1165[31:0];
  _RAND_1166 = {1{`RANDOM}};
  stage4_regs_10_1_4 = _RAND_1166[31:0];
  _RAND_1167 = {1{`RANDOM}};
  stage4_regs_10_1_5 = _RAND_1167[31:0];
  _RAND_1168 = {1{`RANDOM}};
  stage4_regs_10_1_6 = _RAND_1168[31:0];
  _RAND_1169 = {1{`RANDOM}};
  stage4_regs_10_1_7 = _RAND_1169[31:0];
  _RAND_1170 = {1{`RANDOM}};
  stage4_regs_10_1_8 = _RAND_1170[31:0];
  _RAND_1171 = {1{`RANDOM}};
  stage4_regs_11_1_0 = _RAND_1171[31:0];
  _RAND_1172 = {1{`RANDOM}};
  stage4_regs_11_1_1 = _RAND_1172[31:0];
  _RAND_1173 = {1{`RANDOM}};
  stage4_regs_11_1_2 = _RAND_1173[31:0];
  _RAND_1174 = {1{`RANDOM}};
  stage4_regs_11_1_3 = _RAND_1174[31:0];
  _RAND_1175 = {1{`RANDOM}};
  stage4_regs_11_1_4 = _RAND_1175[31:0];
  _RAND_1176 = {1{`RANDOM}};
  stage4_regs_11_1_5 = _RAND_1176[31:0];
  _RAND_1177 = {1{`RANDOM}};
  stage4_regs_11_1_6 = _RAND_1177[31:0];
  _RAND_1178 = {1{`RANDOM}};
  stage4_regs_11_1_7 = _RAND_1178[31:0];
  _RAND_1179 = {1{`RANDOM}};
  stage4_regs_11_1_8 = _RAND_1179[31:0];
  _RAND_1180 = {1{`RANDOM}};
  stage4_regs_12_1_0 = _RAND_1180[31:0];
  _RAND_1181 = {1{`RANDOM}};
  stage4_regs_12_1_1 = _RAND_1181[31:0];
  _RAND_1182 = {1{`RANDOM}};
  stage4_regs_12_1_2 = _RAND_1182[31:0];
  _RAND_1183 = {1{`RANDOM}};
  stage4_regs_12_1_3 = _RAND_1183[31:0];
  _RAND_1184 = {1{`RANDOM}};
  stage4_regs_12_1_4 = _RAND_1184[31:0];
  _RAND_1185 = {1{`RANDOM}};
  stage4_regs_12_1_5 = _RAND_1185[31:0];
  _RAND_1186 = {1{`RANDOM}};
  stage4_regs_12_1_6 = _RAND_1186[31:0];
  _RAND_1187 = {1{`RANDOM}};
  stage4_regs_12_1_7 = _RAND_1187[31:0];
  _RAND_1188 = {1{`RANDOM}};
  stage4_regs_12_1_8 = _RAND_1188[31:0];
  _RAND_1189 = {1{`RANDOM}};
  stage4_regs_13_1_0 = _RAND_1189[31:0];
  _RAND_1190 = {1{`RANDOM}};
  stage4_regs_13_1_1 = _RAND_1190[31:0];
  _RAND_1191 = {1{`RANDOM}};
  stage4_regs_13_1_2 = _RAND_1191[31:0];
  _RAND_1192 = {1{`RANDOM}};
  stage4_regs_13_1_3 = _RAND_1192[31:0];
  _RAND_1193 = {1{`RANDOM}};
  stage4_regs_13_1_4 = _RAND_1193[31:0];
  _RAND_1194 = {1{`RANDOM}};
  stage4_regs_13_1_5 = _RAND_1194[31:0];
  _RAND_1195 = {1{`RANDOM}};
  stage4_regs_13_1_6 = _RAND_1195[31:0];
  _RAND_1196 = {1{`RANDOM}};
  stage4_regs_13_1_7 = _RAND_1196[31:0];
  _RAND_1197 = {1{`RANDOM}};
  stage4_regs_13_1_8 = _RAND_1197[31:0];
  _RAND_1198 = {1{`RANDOM}};
  stage4_regs_14_1_0 = _RAND_1198[31:0];
  _RAND_1199 = {1{`RANDOM}};
  stage4_regs_14_1_1 = _RAND_1199[31:0];
  _RAND_1200 = {1{`RANDOM}};
  stage4_regs_14_1_2 = _RAND_1200[31:0];
  _RAND_1201 = {1{`RANDOM}};
  stage4_regs_14_1_3 = _RAND_1201[31:0];
  _RAND_1202 = {1{`RANDOM}};
  stage4_regs_14_1_4 = _RAND_1202[31:0];
  _RAND_1203 = {1{`RANDOM}};
  stage4_regs_14_1_5 = _RAND_1203[31:0];
  _RAND_1204 = {1{`RANDOM}};
  stage4_regs_14_1_6 = _RAND_1204[31:0];
  _RAND_1205 = {1{`RANDOM}};
  stage4_regs_14_1_7 = _RAND_1205[31:0];
  _RAND_1206 = {1{`RANDOM}};
  stage4_regs_14_1_8 = _RAND_1206[31:0];
  _RAND_1207 = {1{`RANDOM}};
  stage4_regs_15_1_0 = _RAND_1207[31:0];
  _RAND_1208 = {1{`RANDOM}};
  stage4_regs_15_1_1 = _RAND_1208[31:0];
  _RAND_1209 = {1{`RANDOM}};
  stage4_regs_15_1_2 = _RAND_1209[31:0];
  _RAND_1210 = {1{`RANDOM}};
  stage4_regs_15_1_3 = _RAND_1210[31:0];
  _RAND_1211 = {1{`RANDOM}};
  stage4_regs_15_1_4 = _RAND_1211[31:0];
  _RAND_1212 = {1{`RANDOM}};
  stage4_regs_15_1_5 = _RAND_1212[31:0];
  _RAND_1213 = {1{`RANDOM}};
  stage4_regs_15_1_6 = _RAND_1213[31:0];
  _RAND_1214 = {1{`RANDOM}};
  stage4_regs_15_1_7 = _RAND_1214[31:0];
  _RAND_1215 = {1{`RANDOM}};
  stage4_regs_15_1_8 = _RAND_1215[31:0];
  _RAND_1216 = {1{`RANDOM}};
  a_2_isr_to_r = _RAND_1216[31:0];
  _RAND_1217 = {1{`RANDOM}};
  transition_regs_0 = _RAND_1217[31:0];
  _RAND_1218 = {1{`RANDOM}};
  transition_regs_1 = _RAND_1218[31:0];
  _RAND_1219 = {1{`RANDOM}};
  transition_regs_2 = _RAND_1219[31:0];
  _RAND_1220 = {1{`RANDOM}};
  transition_regs_3 = _RAND_1220[31:0];
  _RAND_1221 = {1{`RANDOM}};
  transition_regs_4 = _RAND_1221[31:0];
  _RAND_1222 = {1{`RANDOM}};
  transition_regs_5 = _RAND_1222[31:0];
  _RAND_1223 = {1{`RANDOM}};
  transition_regs_6 = _RAND_1223[31:0];
  _RAND_1224 = {1{`RANDOM}};
  transition_regs_7 = _RAND_1224[31:0];
  _RAND_1225 = {1{`RANDOM}};
  transition_regs_8 = _RAND_1225[31:0];
  _RAND_1226 = {1{`RANDOM}};
  x_n_r_0 = _RAND_1226[31:0];
  _RAND_1227 = {1{`RANDOM}};
  x_n_r_1 = _RAND_1227[31:0];
  _RAND_1228 = {1{`RANDOM}};
  x_n_r_3 = _RAND_1228[31:0];
  _RAND_1229 = {1{`RANDOM}};
  x_n_r_4 = _RAND_1229[31:0];
  _RAND_1230 = {1{`RANDOM}};
  x_n_r_6 = _RAND_1230[31:0];
  _RAND_1231 = {1{`RANDOM}};
  x_n_r_7 = _RAND_1231[31:0];
  _RAND_1232 = {1{`RANDOM}};
  x_n_r_9 = _RAND_1232[31:0];
  _RAND_1233 = {1{`RANDOM}};
  x_n_r_10 = _RAND_1233[31:0];
  _RAND_1234 = {1{`RANDOM}};
  x_n_r_12 = _RAND_1234[31:0];
  _RAND_1235 = {1{`RANDOM}};
  x_n_r_13 = _RAND_1235[31:0];
  _RAND_1236 = {1{`RANDOM}};
  x_n_r_15 = _RAND_1236[31:0];
  _RAND_1237 = {1{`RANDOM}};
  x_n_r_16 = _RAND_1237[31:0];
  _RAND_1238 = {1{`RANDOM}};
  x_n_r_18 = _RAND_1238[31:0];
  _RAND_1239 = {1{`RANDOM}};
  x_n_r_19 = _RAND_1239[31:0];
  _RAND_1240 = {1{`RANDOM}};
  x_n_r_21 = _RAND_1240[31:0];
  _RAND_1241 = {1{`RANDOM}};
  x_n_r_22 = _RAND_1241[31:0];
  _RAND_1242 = {1{`RANDOM}};
  x_n_r_24 = _RAND_1242[31:0];
  _RAND_1243 = {1{`RANDOM}};
  x_n_r_25 = _RAND_1243[31:0];
  _RAND_1244 = {1{`RANDOM}};
  x_n_r_27 = _RAND_1244[31:0];
  _RAND_1245 = {1{`RANDOM}};
  x_n_r_28 = _RAND_1245[31:0];
  _RAND_1246 = {1{`RANDOM}};
  x_n_r_30 = _RAND_1246[31:0];
  _RAND_1247 = {1{`RANDOM}};
  x_n_r_31 = _RAND_1247[31:0];
  _RAND_1248 = {1{`RANDOM}};
  x_n_r_33 = _RAND_1248[31:0];
  _RAND_1249 = {1{`RANDOM}};
  x_n_r_34 = _RAND_1249[31:0];
  _RAND_1250 = {1{`RANDOM}};
  x_n_r_36 = _RAND_1250[31:0];
  _RAND_1251 = {1{`RANDOM}};
  x_n_r_37 = _RAND_1251[31:0];
  _RAND_1252 = {1{`RANDOM}};
  x_n_r_39 = _RAND_1252[31:0];
  _RAND_1253 = {1{`RANDOM}};
  x_n_r_40 = _RAND_1253[31:0];
  _RAND_1254 = {1{`RANDOM}};
  x_n_r_42 = _RAND_1254[31:0];
  _RAND_1255 = {1{`RANDOM}};
  x_n_r_43 = _RAND_1255[31:0];
  _RAND_1256 = {1{`RANDOM}};
  x_n_r_45 = _RAND_1256[31:0];
  _RAND_1257 = {1{`RANDOM}};
  x_n_r_46 = _RAND_1257[31:0];
  _RAND_1258 = {1{`RANDOM}};
  x_n_r_48 = _RAND_1258[31:0];
  _RAND_1259 = {1{`RANDOM}};
  x_n_r_49 = _RAND_1259[31:0];
  _RAND_1260 = {1{`RANDOM}};
  a_2_r_0 = _RAND_1260[31:0];
  _RAND_1261 = {1{`RANDOM}};
  a_2_r_1 = _RAND_1261[31:0];
  _RAND_1262 = {1{`RANDOM}};
  a_2_r_2 = _RAND_1262[31:0];
  _RAND_1263 = {1{`RANDOM}};
  a_2_r_3 = _RAND_1263[31:0];
  _RAND_1264 = {1{`RANDOM}};
  a_2_r_4 = _RAND_1264[31:0];
  _RAND_1265 = {1{`RANDOM}};
  a_2_r_5 = _RAND_1265[31:0];
  _RAND_1266 = {1{`RANDOM}};
  a_2_r_6 = _RAND_1266[31:0];
  _RAND_1267 = {1{`RANDOM}};
  a_2_r_7 = _RAND_1267[31:0];
  _RAND_1268 = {1{`RANDOM}};
  a_2_r_8 = _RAND_1268[31:0];
  _RAND_1269 = {1{`RANDOM}};
  a_2_r_9 = _RAND_1269[31:0];
  _RAND_1270 = {1{`RANDOM}};
  a_2_r_10 = _RAND_1270[31:0];
  _RAND_1271 = {1{`RANDOM}};
  a_2_r_11 = _RAND_1271[31:0];
  _RAND_1272 = {1{`RANDOM}};
  a_2_r_12 = _RAND_1272[31:0];
  _RAND_1273 = {1{`RANDOM}};
  a_2_r_13 = _RAND_1273[31:0];
  _RAND_1274 = {1{`RANDOM}};
  a_2_r_14 = _RAND_1274[31:0];
  _RAND_1275 = {1{`RANDOM}};
  a_2_r_15 = _RAND_1275[31:0];
  _RAND_1276 = {1{`RANDOM}};
  a_2_r_16 = _RAND_1276[31:0];
  _RAND_1277 = {1{`RANDOM}};
  a_2_r_17 = _RAND_1277[31:0];
  _RAND_1278 = {1{`RANDOM}};
  a_2_r_18 = _RAND_1278[31:0];
  _RAND_1279 = {1{`RANDOM}};
  a_2_r_19 = _RAND_1279[31:0];
  _RAND_1280 = {1{`RANDOM}};
  a_2_r_20 = _RAND_1280[31:0];
  _RAND_1281 = {1{`RANDOM}};
  a_2_r_21 = _RAND_1281[31:0];
  _RAND_1282 = {1{`RANDOM}};
  a_2_r_22 = _RAND_1282[31:0];
  _RAND_1283 = {1{`RANDOM}};
  a_2_r_23 = _RAND_1283[31:0];
  _RAND_1284 = {1{`RANDOM}};
  a_2_r_24 = _RAND_1284[31:0];
  _RAND_1285 = {1{`RANDOM}};
  a_2_r_25 = _RAND_1285[31:0];
  _RAND_1286 = {1{`RANDOM}};
  a_2_r_26 = _RAND_1286[31:0];
  _RAND_1287 = {1{`RANDOM}};
  a_2_r_27 = _RAND_1287[31:0];
  _RAND_1288 = {1{`RANDOM}};
  a_2_r_28 = _RAND_1288[31:0];
  _RAND_1289 = {1{`RANDOM}};
  a_2_r_29 = _RAND_1289[31:0];
  _RAND_1290 = {1{`RANDOM}};
  a_2_r_30 = _RAND_1290[31:0];
  _RAND_1291 = {1{`RANDOM}};
  a_2_r_31 = _RAND_1291[31:0];
  _RAND_1292 = {1{`RANDOM}};
  a_2_r_32 = _RAND_1292[31:0];
  _RAND_1293 = {1{`RANDOM}};
  a_2_r_33 = _RAND_1293[31:0];
  _RAND_1294 = {1{`RANDOM}};
  a_2_r_34 = _RAND_1294[31:0];
  _RAND_1295 = {1{`RANDOM}};
  a_2_r_35 = _RAND_1295[31:0];
  _RAND_1296 = {1{`RANDOM}};
  a_2_r_36 = _RAND_1296[31:0];
  _RAND_1297 = {1{`RANDOM}};
  a_2_r_37 = _RAND_1297[31:0];
  _RAND_1298 = {1{`RANDOM}};
  a_2_r_38 = _RAND_1298[31:0];
  _RAND_1299 = {1{`RANDOM}};
  a_2_r_39 = _RAND_1299[31:0];
  _RAND_1300 = {1{`RANDOM}};
  a_2_r_40 = _RAND_1300[31:0];
  _RAND_1301 = {1{`RANDOM}};
  a_2_r_41 = _RAND_1301[31:0];
  _RAND_1302 = {1{`RANDOM}};
  a_2_r_42 = _RAND_1302[31:0];
  _RAND_1303 = {1{`RANDOM}};
  a_2_r_43 = _RAND_1303[31:0];
  _RAND_1304 = {1{`RANDOM}};
  a_2_r_44 = _RAND_1304[31:0];
  _RAND_1305 = {1{`RANDOM}};
  a_2_r_45 = _RAND_1305[31:0];
  _RAND_1306 = {1{`RANDOM}};
  a_2_r_46 = _RAND_1306[31:0];
  _RAND_1307 = {1{`RANDOM}};
  a_2_r_47 = _RAND_1307[31:0];
  _RAND_1308 = {1{`RANDOM}};
  a_2_r_48 = _RAND_1308[31:0];
  _RAND_1309 = {1{`RANDOM}};
  a_2_r_49 = _RAND_1309[31:0];
  _RAND_1310 = {1{`RANDOM}};
  a_2_r_50 = _RAND_1310[31:0];
  _RAND_1311 = {1{`RANDOM}};
  stage1_regs_r_0_0_0 = _RAND_1311[31:0];
  _RAND_1312 = {1{`RANDOM}};
  stage1_regs_r_0_0_1 = _RAND_1312[31:0];
  _RAND_1313 = {1{`RANDOM}};
  stage1_regs_r_0_0_2 = _RAND_1313[31:0];
  _RAND_1314 = {1{`RANDOM}};
  stage1_regs_r_0_0_3 = _RAND_1314[31:0];
  _RAND_1315 = {1{`RANDOM}};
  stage1_regs_r_0_0_4 = _RAND_1315[31:0];
  _RAND_1316 = {1{`RANDOM}};
  stage1_regs_r_0_0_5 = _RAND_1316[31:0];
  _RAND_1317 = {1{`RANDOM}};
  stage1_regs_r_0_0_6 = _RAND_1317[31:0];
  _RAND_1318 = {1{`RANDOM}};
  stage1_regs_r_0_0_7 = _RAND_1318[31:0];
  _RAND_1319 = {1{`RANDOM}};
  stage1_regs_r_0_0_8 = _RAND_1319[31:0];
  _RAND_1320 = {1{`RANDOM}};
  stage1_regs_r_0_1_0 = _RAND_1320[31:0];
  _RAND_1321 = {1{`RANDOM}};
  stage1_regs_r_0_1_1 = _RAND_1321[31:0];
  _RAND_1322 = {1{`RANDOM}};
  stage1_regs_r_0_1_2 = _RAND_1322[31:0];
  _RAND_1323 = {1{`RANDOM}};
  stage1_regs_r_0_1_3 = _RAND_1323[31:0];
  _RAND_1324 = {1{`RANDOM}};
  stage1_regs_r_0_1_4 = _RAND_1324[31:0];
  _RAND_1325 = {1{`RANDOM}};
  stage1_regs_r_0_1_5 = _RAND_1325[31:0];
  _RAND_1326 = {1{`RANDOM}};
  stage1_regs_r_0_1_6 = _RAND_1326[31:0];
  _RAND_1327 = {1{`RANDOM}};
  stage1_regs_r_0_1_7 = _RAND_1327[31:0];
  _RAND_1328 = {1{`RANDOM}};
  stage1_regs_r_0_1_8 = _RAND_1328[31:0];
  _RAND_1329 = {1{`RANDOM}};
  stage1_regs_r_1_0_0 = _RAND_1329[31:0];
  _RAND_1330 = {1{`RANDOM}};
  stage1_regs_r_1_0_1 = _RAND_1330[31:0];
  _RAND_1331 = {1{`RANDOM}};
  stage1_regs_r_1_0_2 = _RAND_1331[31:0];
  _RAND_1332 = {1{`RANDOM}};
  stage1_regs_r_1_0_3 = _RAND_1332[31:0];
  _RAND_1333 = {1{`RANDOM}};
  stage1_regs_r_1_0_4 = _RAND_1333[31:0];
  _RAND_1334 = {1{`RANDOM}};
  stage1_regs_r_1_0_5 = _RAND_1334[31:0];
  _RAND_1335 = {1{`RANDOM}};
  stage1_regs_r_1_0_6 = _RAND_1335[31:0];
  _RAND_1336 = {1{`RANDOM}};
  stage1_regs_r_1_0_7 = _RAND_1336[31:0];
  _RAND_1337 = {1{`RANDOM}};
  stage1_regs_r_1_0_8 = _RAND_1337[31:0];
  _RAND_1338 = {1{`RANDOM}};
  stage1_regs_r_1_1_0 = _RAND_1338[31:0];
  _RAND_1339 = {1{`RANDOM}};
  stage1_regs_r_1_1_1 = _RAND_1339[31:0];
  _RAND_1340 = {1{`RANDOM}};
  stage1_regs_r_1_1_2 = _RAND_1340[31:0];
  _RAND_1341 = {1{`RANDOM}};
  stage1_regs_r_1_1_3 = _RAND_1341[31:0];
  _RAND_1342 = {1{`RANDOM}};
  stage1_regs_r_1_1_4 = _RAND_1342[31:0];
  _RAND_1343 = {1{`RANDOM}};
  stage1_regs_r_1_1_5 = _RAND_1343[31:0];
  _RAND_1344 = {1{`RANDOM}};
  stage1_regs_r_1_1_6 = _RAND_1344[31:0];
  _RAND_1345 = {1{`RANDOM}};
  stage1_regs_r_1_1_7 = _RAND_1345[31:0];
  _RAND_1346 = {1{`RANDOM}};
  stage1_regs_r_1_1_8 = _RAND_1346[31:0];
  _RAND_1347 = {1{`RANDOM}};
  stage1_regs_r_2_0_0 = _RAND_1347[31:0];
  _RAND_1348 = {1{`RANDOM}};
  stage1_regs_r_2_0_1 = _RAND_1348[31:0];
  _RAND_1349 = {1{`RANDOM}};
  stage1_regs_r_2_0_2 = _RAND_1349[31:0];
  _RAND_1350 = {1{`RANDOM}};
  stage1_regs_r_2_0_3 = _RAND_1350[31:0];
  _RAND_1351 = {1{`RANDOM}};
  stage1_regs_r_2_0_4 = _RAND_1351[31:0];
  _RAND_1352 = {1{`RANDOM}};
  stage1_regs_r_2_0_5 = _RAND_1352[31:0];
  _RAND_1353 = {1{`RANDOM}};
  stage1_regs_r_2_0_6 = _RAND_1353[31:0];
  _RAND_1354 = {1{`RANDOM}};
  stage1_regs_r_2_0_7 = _RAND_1354[31:0];
  _RAND_1355 = {1{`RANDOM}};
  stage1_regs_r_2_0_8 = _RAND_1355[31:0];
  _RAND_1356 = {1{`RANDOM}};
  stage1_regs_r_2_1_0 = _RAND_1356[31:0];
  _RAND_1357 = {1{`RANDOM}};
  stage1_regs_r_2_1_1 = _RAND_1357[31:0];
  _RAND_1358 = {1{`RANDOM}};
  stage1_regs_r_2_1_2 = _RAND_1358[31:0];
  _RAND_1359 = {1{`RANDOM}};
  stage1_regs_r_2_1_3 = _RAND_1359[31:0];
  _RAND_1360 = {1{`RANDOM}};
  stage1_regs_r_2_1_4 = _RAND_1360[31:0];
  _RAND_1361 = {1{`RANDOM}};
  stage1_regs_r_2_1_5 = _RAND_1361[31:0];
  _RAND_1362 = {1{`RANDOM}};
  stage1_regs_r_2_1_6 = _RAND_1362[31:0];
  _RAND_1363 = {1{`RANDOM}};
  stage1_regs_r_2_1_7 = _RAND_1363[31:0];
  _RAND_1364 = {1{`RANDOM}};
  stage1_regs_r_2_1_8 = _RAND_1364[31:0];
  _RAND_1365 = {1{`RANDOM}};
  stage1_regs_r_3_0_0 = _RAND_1365[31:0];
  _RAND_1366 = {1{`RANDOM}};
  stage1_regs_r_3_0_1 = _RAND_1366[31:0];
  _RAND_1367 = {1{`RANDOM}};
  stage1_regs_r_3_0_2 = _RAND_1367[31:0];
  _RAND_1368 = {1{`RANDOM}};
  stage1_regs_r_3_0_3 = _RAND_1368[31:0];
  _RAND_1369 = {1{`RANDOM}};
  stage1_regs_r_3_0_4 = _RAND_1369[31:0];
  _RAND_1370 = {1{`RANDOM}};
  stage1_regs_r_3_0_5 = _RAND_1370[31:0];
  _RAND_1371 = {1{`RANDOM}};
  stage1_regs_r_3_0_6 = _RAND_1371[31:0];
  _RAND_1372 = {1{`RANDOM}};
  stage1_regs_r_3_0_7 = _RAND_1372[31:0];
  _RAND_1373 = {1{`RANDOM}};
  stage1_regs_r_3_0_8 = _RAND_1373[31:0];
  _RAND_1374 = {1{`RANDOM}};
  stage1_regs_r_3_1_0 = _RAND_1374[31:0];
  _RAND_1375 = {1{`RANDOM}};
  stage1_regs_r_3_1_1 = _RAND_1375[31:0];
  _RAND_1376 = {1{`RANDOM}};
  stage1_regs_r_3_1_2 = _RAND_1376[31:0];
  _RAND_1377 = {1{`RANDOM}};
  stage1_regs_r_3_1_3 = _RAND_1377[31:0];
  _RAND_1378 = {1{`RANDOM}};
  stage1_regs_r_3_1_4 = _RAND_1378[31:0];
  _RAND_1379 = {1{`RANDOM}};
  stage1_regs_r_3_1_5 = _RAND_1379[31:0];
  _RAND_1380 = {1{`RANDOM}};
  stage1_regs_r_3_1_6 = _RAND_1380[31:0];
  _RAND_1381 = {1{`RANDOM}};
  stage1_regs_r_3_1_7 = _RAND_1381[31:0];
  _RAND_1382 = {1{`RANDOM}};
  stage1_regs_r_3_1_8 = _RAND_1382[31:0];
  _RAND_1383 = {1{`RANDOM}};
  stage1_regs_r_4_0_0 = _RAND_1383[31:0];
  _RAND_1384 = {1{`RANDOM}};
  stage1_regs_r_4_0_1 = _RAND_1384[31:0];
  _RAND_1385 = {1{`RANDOM}};
  stage1_regs_r_4_0_2 = _RAND_1385[31:0];
  _RAND_1386 = {1{`RANDOM}};
  stage1_regs_r_4_0_3 = _RAND_1386[31:0];
  _RAND_1387 = {1{`RANDOM}};
  stage1_regs_r_4_0_4 = _RAND_1387[31:0];
  _RAND_1388 = {1{`RANDOM}};
  stage1_regs_r_4_0_5 = _RAND_1388[31:0];
  _RAND_1389 = {1{`RANDOM}};
  stage1_regs_r_4_0_6 = _RAND_1389[31:0];
  _RAND_1390 = {1{`RANDOM}};
  stage1_regs_r_4_0_7 = _RAND_1390[31:0];
  _RAND_1391 = {1{`RANDOM}};
  stage1_regs_r_4_0_8 = _RAND_1391[31:0];
  _RAND_1392 = {1{`RANDOM}};
  stage1_regs_r_4_1_0 = _RAND_1392[31:0];
  _RAND_1393 = {1{`RANDOM}};
  stage1_regs_r_4_1_1 = _RAND_1393[31:0];
  _RAND_1394 = {1{`RANDOM}};
  stage1_regs_r_4_1_2 = _RAND_1394[31:0];
  _RAND_1395 = {1{`RANDOM}};
  stage1_regs_r_4_1_3 = _RAND_1395[31:0];
  _RAND_1396 = {1{`RANDOM}};
  stage1_regs_r_4_1_4 = _RAND_1396[31:0];
  _RAND_1397 = {1{`RANDOM}};
  stage1_regs_r_4_1_5 = _RAND_1397[31:0];
  _RAND_1398 = {1{`RANDOM}};
  stage1_regs_r_4_1_6 = _RAND_1398[31:0];
  _RAND_1399 = {1{`RANDOM}};
  stage1_regs_r_4_1_7 = _RAND_1399[31:0];
  _RAND_1400 = {1{`RANDOM}};
  stage1_regs_r_4_1_8 = _RAND_1400[31:0];
  _RAND_1401 = {1{`RANDOM}};
  stage1_regs_r_5_0_0 = _RAND_1401[31:0];
  _RAND_1402 = {1{`RANDOM}};
  stage1_regs_r_5_0_1 = _RAND_1402[31:0];
  _RAND_1403 = {1{`RANDOM}};
  stage1_regs_r_5_0_2 = _RAND_1403[31:0];
  _RAND_1404 = {1{`RANDOM}};
  stage1_regs_r_5_0_3 = _RAND_1404[31:0];
  _RAND_1405 = {1{`RANDOM}};
  stage1_regs_r_5_0_4 = _RAND_1405[31:0];
  _RAND_1406 = {1{`RANDOM}};
  stage1_regs_r_5_0_5 = _RAND_1406[31:0];
  _RAND_1407 = {1{`RANDOM}};
  stage1_regs_r_5_0_6 = _RAND_1407[31:0];
  _RAND_1408 = {1{`RANDOM}};
  stage1_regs_r_5_0_7 = _RAND_1408[31:0];
  _RAND_1409 = {1{`RANDOM}};
  stage1_regs_r_5_0_8 = _RAND_1409[31:0];
  _RAND_1410 = {1{`RANDOM}};
  stage1_regs_r_5_1_0 = _RAND_1410[31:0];
  _RAND_1411 = {1{`RANDOM}};
  stage1_regs_r_5_1_1 = _RAND_1411[31:0];
  _RAND_1412 = {1{`RANDOM}};
  stage1_regs_r_5_1_2 = _RAND_1412[31:0];
  _RAND_1413 = {1{`RANDOM}};
  stage1_regs_r_5_1_3 = _RAND_1413[31:0];
  _RAND_1414 = {1{`RANDOM}};
  stage1_regs_r_5_1_4 = _RAND_1414[31:0];
  _RAND_1415 = {1{`RANDOM}};
  stage1_regs_r_5_1_5 = _RAND_1415[31:0];
  _RAND_1416 = {1{`RANDOM}};
  stage1_regs_r_5_1_6 = _RAND_1416[31:0];
  _RAND_1417 = {1{`RANDOM}};
  stage1_regs_r_5_1_7 = _RAND_1417[31:0];
  _RAND_1418 = {1{`RANDOM}};
  stage1_regs_r_5_1_8 = _RAND_1418[31:0];
  _RAND_1419 = {1{`RANDOM}};
  stage1_regs_r_6_0_0 = _RAND_1419[31:0];
  _RAND_1420 = {1{`RANDOM}};
  stage1_regs_r_6_0_1 = _RAND_1420[31:0];
  _RAND_1421 = {1{`RANDOM}};
  stage1_regs_r_6_0_2 = _RAND_1421[31:0];
  _RAND_1422 = {1{`RANDOM}};
  stage1_regs_r_6_0_3 = _RAND_1422[31:0];
  _RAND_1423 = {1{`RANDOM}};
  stage1_regs_r_6_0_4 = _RAND_1423[31:0];
  _RAND_1424 = {1{`RANDOM}};
  stage1_regs_r_6_0_5 = _RAND_1424[31:0];
  _RAND_1425 = {1{`RANDOM}};
  stage1_regs_r_6_0_6 = _RAND_1425[31:0];
  _RAND_1426 = {1{`RANDOM}};
  stage1_regs_r_6_0_7 = _RAND_1426[31:0];
  _RAND_1427 = {1{`RANDOM}};
  stage1_regs_r_6_0_8 = _RAND_1427[31:0];
  _RAND_1428 = {1{`RANDOM}};
  stage1_regs_r_6_1_0 = _RAND_1428[31:0];
  _RAND_1429 = {1{`RANDOM}};
  stage1_regs_r_6_1_1 = _RAND_1429[31:0];
  _RAND_1430 = {1{`RANDOM}};
  stage1_regs_r_6_1_2 = _RAND_1430[31:0];
  _RAND_1431 = {1{`RANDOM}};
  stage1_regs_r_6_1_3 = _RAND_1431[31:0];
  _RAND_1432 = {1{`RANDOM}};
  stage1_regs_r_6_1_4 = _RAND_1432[31:0];
  _RAND_1433 = {1{`RANDOM}};
  stage1_regs_r_6_1_5 = _RAND_1433[31:0];
  _RAND_1434 = {1{`RANDOM}};
  stage1_regs_r_6_1_6 = _RAND_1434[31:0];
  _RAND_1435 = {1{`RANDOM}};
  stage1_regs_r_6_1_7 = _RAND_1435[31:0];
  _RAND_1436 = {1{`RANDOM}};
  stage1_regs_r_6_1_8 = _RAND_1436[31:0];
  _RAND_1437 = {1{`RANDOM}};
  stage1_regs_r_7_0_0 = _RAND_1437[31:0];
  _RAND_1438 = {1{`RANDOM}};
  stage1_regs_r_7_0_1 = _RAND_1438[31:0];
  _RAND_1439 = {1{`RANDOM}};
  stage1_regs_r_7_0_2 = _RAND_1439[31:0];
  _RAND_1440 = {1{`RANDOM}};
  stage1_regs_r_7_0_3 = _RAND_1440[31:0];
  _RAND_1441 = {1{`RANDOM}};
  stage1_regs_r_7_0_4 = _RAND_1441[31:0];
  _RAND_1442 = {1{`RANDOM}};
  stage1_regs_r_7_0_5 = _RAND_1442[31:0];
  _RAND_1443 = {1{`RANDOM}};
  stage1_regs_r_7_0_6 = _RAND_1443[31:0];
  _RAND_1444 = {1{`RANDOM}};
  stage1_regs_r_7_0_7 = _RAND_1444[31:0];
  _RAND_1445 = {1{`RANDOM}};
  stage1_regs_r_7_0_8 = _RAND_1445[31:0];
  _RAND_1446 = {1{`RANDOM}};
  stage1_regs_r_7_1_0 = _RAND_1446[31:0];
  _RAND_1447 = {1{`RANDOM}};
  stage1_regs_r_7_1_1 = _RAND_1447[31:0];
  _RAND_1448 = {1{`RANDOM}};
  stage1_regs_r_7_1_2 = _RAND_1448[31:0];
  _RAND_1449 = {1{`RANDOM}};
  stage1_regs_r_7_1_3 = _RAND_1449[31:0];
  _RAND_1450 = {1{`RANDOM}};
  stage1_regs_r_7_1_4 = _RAND_1450[31:0];
  _RAND_1451 = {1{`RANDOM}};
  stage1_regs_r_7_1_5 = _RAND_1451[31:0];
  _RAND_1452 = {1{`RANDOM}};
  stage1_regs_r_7_1_6 = _RAND_1452[31:0];
  _RAND_1453 = {1{`RANDOM}};
  stage1_regs_r_7_1_7 = _RAND_1453[31:0];
  _RAND_1454 = {1{`RANDOM}};
  stage1_regs_r_7_1_8 = _RAND_1454[31:0];
  _RAND_1455 = {1{`RANDOM}};
  stage1_regs_r_8_0_0 = _RAND_1455[31:0];
  _RAND_1456 = {1{`RANDOM}};
  stage1_regs_r_8_0_1 = _RAND_1456[31:0];
  _RAND_1457 = {1{`RANDOM}};
  stage1_regs_r_8_0_2 = _RAND_1457[31:0];
  _RAND_1458 = {1{`RANDOM}};
  stage1_regs_r_8_0_3 = _RAND_1458[31:0];
  _RAND_1459 = {1{`RANDOM}};
  stage1_regs_r_8_0_4 = _RAND_1459[31:0];
  _RAND_1460 = {1{`RANDOM}};
  stage1_regs_r_8_0_5 = _RAND_1460[31:0];
  _RAND_1461 = {1{`RANDOM}};
  stage1_regs_r_8_0_6 = _RAND_1461[31:0];
  _RAND_1462 = {1{`RANDOM}};
  stage1_regs_r_8_0_7 = _RAND_1462[31:0];
  _RAND_1463 = {1{`RANDOM}};
  stage1_regs_r_8_0_8 = _RAND_1463[31:0];
  _RAND_1464 = {1{`RANDOM}};
  stage1_regs_r_8_1_0 = _RAND_1464[31:0];
  _RAND_1465 = {1{`RANDOM}};
  stage1_regs_r_8_1_1 = _RAND_1465[31:0];
  _RAND_1466 = {1{`RANDOM}};
  stage1_regs_r_8_1_2 = _RAND_1466[31:0];
  _RAND_1467 = {1{`RANDOM}};
  stage1_regs_r_8_1_3 = _RAND_1467[31:0];
  _RAND_1468 = {1{`RANDOM}};
  stage1_regs_r_8_1_4 = _RAND_1468[31:0];
  _RAND_1469 = {1{`RANDOM}};
  stage1_regs_r_8_1_5 = _RAND_1469[31:0];
  _RAND_1470 = {1{`RANDOM}};
  stage1_regs_r_8_1_6 = _RAND_1470[31:0];
  _RAND_1471 = {1{`RANDOM}};
  stage1_regs_r_8_1_7 = _RAND_1471[31:0];
  _RAND_1472 = {1{`RANDOM}};
  stage1_regs_r_8_1_8 = _RAND_1472[31:0];
  _RAND_1473 = {1{`RANDOM}};
  stage1_regs_r_9_0_0 = _RAND_1473[31:0];
  _RAND_1474 = {1{`RANDOM}};
  stage1_regs_r_9_0_1 = _RAND_1474[31:0];
  _RAND_1475 = {1{`RANDOM}};
  stage1_regs_r_9_0_2 = _RAND_1475[31:0];
  _RAND_1476 = {1{`RANDOM}};
  stage1_regs_r_9_0_3 = _RAND_1476[31:0];
  _RAND_1477 = {1{`RANDOM}};
  stage1_regs_r_9_0_4 = _RAND_1477[31:0];
  _RAND_1478 = {1{`RANDOM}};
  stage1_regs_r_9_0_5 = _RAND_1478[31:0];
  _RAND_1479 = {1{`RANDOM}};
  stage1_regs_r_9_0_6 = _RAND_1479[31:0];
  _RAND_1480 = {1{`RANDOM}};
  stage1_regs_r_9_0_7 = _RAND_1480[31:0];
  _RAND_1481 = {1{`RANDOM}};
  stage1_regs_r_9_0_8 = _RAND_1481[31:0];
  _RAND_1482 = {1{`RANDOM}};
  stage1_regs_r_9_1_0 = _RAND_1482[31:0];
  _RAND_1483 = {1{`RANDOM}};
  stage1_regs_r_9_1_1 = _RAND_1483[31:0];
  _RAND_1484 = {1{`RANDOM}};
  stage1_regs_r_9_1_2 = _RAND_1484[31:0];
  _RAND_1485 = {1{`RANDOM}};
  stage1_regs_r_9_1_3 = _RAND_1485[31:0];
  _RAND_1486 = {1{`RANDOM}};
  stage1_regs_r_9_1_4 = _RAND_1486[31:0];
  _RAND_1487 = {1{`RANDOM}};
  stage1_regs_r_9_1_5 = _RAND_1487[31:0];
  _RAND_1488 = {1{`RANDOM}};
  stage1_regs_r_9_1_6 = _RAND_1488[31:0];
  _RAND_1489 = {1{`RANDOM}};
  stage1_regs_r_9_1_7 = _RAND_1489[31:0];
  _RAND_1490 = {1{`RANDOM}};
  stage1_regs_r_9_1_8 = _RAND_1490[31:0];
  _RAND_1491 = {1{`RANDOM}};
  stage1_regs_r_10_0_0 = _RAND_1491[31:0];
  _RAND_1492 = {1{`RANDOM}};
  stage1_regs_r_10_0_1 = _RAND_1492[31:0];
  _RAND_1493 = {1{`RANDOM}};
  stage1_regs_r_10_0_2 = _RAND_1493[31:0];
  _RAND_1494 = {1{`RANDOM}};
  stage1_regs_r_10_0_3 = _RAND_1494[31:0];
  _RAND_1495 = {1{`RANDOM}};
  stage1_regs_r_10_0_4 = _RAND_1495[31:0];
  _RAND_1496 = {1{`RANDOM}};
  stage1_regs_r_10_0_5 = _RAND_1496[31:0];
  _RAND_1497 = {1{`RANDOM}};
  stage1_regs_r_10_0_6 = _RAND_1497[31:0];
  _RAND_1498 = {1{`RANDOM}};
  stage1_regs_r_10_0_7 = _RAND_1498[31:0];
  _RAND_1499 = {1{`RANDOM}};
  stage1_regs_r_10_0_8 = _RAND_1499[31:0];
  _RAND_1500 = {1{`RANDOM}};
  stage1_regs_r_10_1_0 = _RAND_1500[31:0];
  _RAND_1501 = {1{`RANDOM}};
  stage1_regs_r_10_1_1 = _RAND_1501[31:0];
  _RAND_1502 = {1{`RANDOM}};
  stage1_regs_r_10_1_2 = _RAND_1502[31:0];
  _RAND_1503 = {1{`RANDOM}};
  stage1_regs_r_10_1_3 = _RAND_1503[31:0];
  _RAND_1504 = {1{`RANDOM}};
  stage1_regs_r_10_1_4 = _RAND_1504[31:0];
  _RAND_1505 = {1{`RANDOM}};
  stage1_regs_r_10_1_5 = _RAND_1505[31:0];
  _RAND_1506 = {1{`RANDOM}};
  stage1_regs_r_10_1_6 = _RAND_1506[31:0];
  _RAND_1507 = {1{`RANDOM}};
  stage1_regs_r_10_1_7 = _RAND_1507[31:0];
  _RAND_1508 = {1{`RANDOM}};
  stage1_regs_r_10_1_8 = _RAND_1508[31:0];
  _RAND_1509 = {1{`RANDOM}};
  stage1_regs_r_11_0_0 = _RAND_1509[31:0];
  _RAND_1510 = {1{`RANDOM}};
  stage1_regs_r_11_0_1 = _RAND_1510[31:0];
  _RAND_1511 = {1{`RANDOM}};
  stage1_regs_r_11_0_2 = _RAND_1511[31:0];
  _RAND_1512 = {1{`RANDOM}};
  stage1_regs_r_11_0_3 = _RAND_1512[31:0];
  _RAND_1513 = {1{`RANDOM}};
  stage1_regs_r_11_0_4 = _RAND_1513[31:0];
  _RAND_1514 = {1{`RANDOM}};
  stage1_regs_r_11_0_5 = _RAND_1514[31:0];
  _RAND_1515 = {1{`RANDOM}};
  stage1_regs_r_11_0_6 = _RAND_1515[31:0];
  _RAND_1516 = {1{`RANDOM}};
  stage1_regs_r_11_0_7 = _RAND_1516[31:0];
  _RAND_1517 = {1{`RANDOM}};
  stage1_regs_r_11_0_8 = _RAND_1517[31:0];
  _RAND_1518 = {1{`RANDOM}};
  stage1_regs_r_11_1_0 = _RAND_1518[31:0];
  _RAND_1519 = {1{`RANDOM}};
  stage1_regs_r_11_1_1 = _RAND_1519[31:0];
  _RAND_1520 = {1{`RANDOM}};
  stage1_regs_r_11_1_2 = _RAND_1520[31:0];
  _RAND_1521 = {1{`RANDOM}};
  stage1_regs_r_11_1_3 = _RAND_1521[31:0];
  _RAND_1522 = {1{`RANDOM}};
  stage1_regs_r_11_1_4 = _RAND_1522[31:0];
  _RAND_1523 = {1{`RANDOM}};
  stage1_regs_r_11_1_5 = _RAND_1523[31:0];
  _RAND_1524 = {1{`RANDOM}};
  stage1_regs_r_11_1_6 = _RAND_1524[31:0];
  _RAND_1525 = {1{`RANDOM}};
  stage1_regs_r_11_1_7 = _RAND_1525[31:0];
  _RAND_1526 = {1{`RANDOM}};
  stage1_regs_r_11_1_8 = _RAND_1526[31:0];
  _RAND_1527 = {1{`RANDOM}};
  stage1_regs_r_12_0_0 = _RAND_1527[31:0];
  _RAND_1528 = {1{`RANDOM}};
  stage1_regs_r_12_0_1 = _RAND_1528[31:0];
  _RAND_1529 = {1{`RANDOM}};
  stage1_regs_r_12_0_2 = _RAND_1529[31:0];
  _RAND_1530 = {1{`RANDOM}};
  stage1_regs_r_12_0_3 = _RAND_1530[31:0];
  _RAND_1531 = {1{`RANDOM}};
  stage1_regs_r_12_0_4 = _RAND_1531[31:0];
  _RAND_1532 = {1{`RANDOM}};
  stage1_regs_r_12_0_5 = _RAND_1532[31:0];
  _RAND_1533 = {1{`RANDOM}};
  stage1_regs_r_12_0_6 = _RAND_1533[31:0];
  _RAND_1534 = {1{`RANDOM}};
  stage1_regs_r_12_0_7 = _RAND_1534[31:0];
  _RAND_1535 = {1{`RANDOM}};
  stage1_regs_r_12_0_8 = _RAND_1535[31:0];
  _RAND_1536 = {1{`RANDOM}};
  stage1_regs_r_12_1_0 = _RAND_1536[31:0];
  _RAND_1537 = {1{`RANDOM}};
  stage1_regs_r_12_1_1 = _RAND_1537[31:0];
  _RAND_1538 = {1{`RANDOM}};
  stage1_regs_r_12_1_2 = _RAND_1538[31:0];
  _RAND_1539 = {1{`RANDOM}};
  stage1_regs_r_12_1_3 = _RAND_1539[31:0];
  _RAND_1540 = {1{`RANDOM}};
  stage1_regs_r_12_1_4 = _RAND_1540[31:0];
  _RAND_1541 = {1{`RANDOM}};
  stage1_regs_r_12_1_5 = _RAND_1541[31:0];
  _RAND_1542 = {1{`RANDOM}};
  stage1_regs_r_12_1_6 = _RAND_1542[31:0];
  _RAND_1543 = {1{`RANDOM}};
  stage1_regs_r_12_1_7 = _RAND_1543[31:0];
  _RAND_1544 = {1{`RANDOM}};
  stage1_regs_r_12_1_8 = _RAND_1544[31:0];
  _RAND_1545 = {1{`RANDOM}};
  stage1_regs_r_13_0_0 = _RAND_1545[31:0];
  _RAND_1546 = {1{`RANDOM}};
  stage1_regs_r_13_0_1 = _RAND_1546[31:0];
  _RAND_1547 = {1{`RANDOM}};
  stage1_regs_r_13_0_2 = _RAND_1547[31:0];
  _RAND_1548 = {1{`RANDOM}};
  stage1_regs_r_13_0_3 = _RAND_1548[31:0];
  _RAND_1549 = {1{`RANDOM}};
  stage1_regs_r_13_0_4 = _RAND_1549[31:0];
  _RAND_1550 = {1{`RANDOM}};
  stage1_regs_r_13_0_5 = _RAND_1550[31:0];
  _RAND_1551 = {1{`RANDOM}};
  stage1_regs_r_13_0_6 = _RAND_1551[31:0];
  _RAND_1552 = {1{`RANDOM}};
  stage1_regs_r_13_0_7 = _RAND_1552[31:0];
  _RAND_1553 = {1{`RANDOM}};
  stage1_regs_r_13_0_8 = _RAND_1553[31:0];
  _RAND_1554 = {1{`RANDOM}};
  stage1_regs_r_13_1_0 = _RAND_1554[31:0];
  _RAND_1555 = {1{`RANDOM}};
  stage1_regs_r_13_1_1 = _RAND_1555[31:0];
  _RAND_1556 = {1{`RANDOM}};
  stage1_regs_r_13_1_2 = _RAND_1556[31:0];
  _RAND_1557 = {1{`RANDOM}};
  stage1_regs_r_13_1_3 = _RAND_1557[31:0];
  _RAND_1558 = {1{`RANDOM}};
  stage1_regs_r_13_1_4 = _RAND_1558[31:0];
  _RAND_1559 = {1{`RANDOM}};
  stage1_regs_r_13_1_5 = _RAND_1559[31:0];
  _RAND_1560 = {1{`RANDOM}};
  stage1_regs_r_13_1_6 = _RAND_1560[31:0];
  _RAND_1561 = {1{`RANDOM}};
  stage1_regs_r_13_1_7 = _RAND_1561[31:0];
  _RAND_1562 = {1{`RANDOM}};
  stage1_regs_r_13_1_8 = _RAND_1562[31:0];
  _RAND_1563 = {1{`RANDOM}};
  stage1_regs_r_14_0_0 = _RAND_1563[31:0];
  _RAND_1564 = {1{`RANDOM}};
  stage1_regs_r_14_0_1 = _RAND_1564[31:0];
  _RAND_1565 = {1{`RANDOM}};
  stage1_regs_r_14_0_2 = _RAND_1565[31:0];
  _RAND_1566 = {1{`RANDOM}};
  stage1_regs_r_14_0_3 = _RAND_1566[31:0];
  _RAND_1567 = {1{`RANDOM}};
  stage1_regs_r_14_0_4 = _RAND_1567[31:0];
  _RAND_1568 = {1{`RANDOM}};
  stage1_regs_r_14_0_5 = _RAND_1568[31:0];
  _RAND_1569 = {1{`RANDOM}};
  stage1_regs_r_14_0_6 = _RAND_1569[31:0];
  _RAND_1570 = {1{`RANDOM}};
  stage1_regs_r_14_0_7 = _RAND_1570[31:0];
  _RAND_1571 = {1{`RANDOM}};
  stage1_regs_r_14_0_8 = _RAND_1571[31:0];
  _RAND_1572 = {1{`RANDOM}};
  stage1_regs_r_14_1_0 = _RAND_1572[31:0];
  _RAND_1573 = {1{`RANDOM}};
  stage1_regs_r_14_1_1 = _RAND_1573[31:0];
  _RAND_1574 = {1{`RANDOM}};
  stage1_regs_r_14_1_2 = _RAND_1574[31:0];
  _RAND_1575 = {1{`RANDOM}};
  stage1_regs_r_14_1_3 = _RAND_1575[31:0];
  _RAND_1576 = {1{`RANDOM}};
  stage1_regs_r_14_1_4 = _RAND_1576[31:0];
  _RAND_1577 = {1{`RANDOM}};
  stage1_regs_r_14_1_5 = _RAND_1577[31:0];
  _RAND_1578 = {1{`RANDOM}};
  stage1_regs_r_14_1_6 = _RAND_1578[31:0];
  _RAND_1579 = {1{`RANDOM}};
  stage1_regs_r_14_1_7 = _RAND_1579[31:0];
  _RAND_1580 = {1{`RANDOM}};
  stage1_regs_r_14_1_8 = _RAND_1580[31:0];
  _RAND_1581 = {1{`RANDOM}};
  stage1_regs_r_15_0_0 = _RAND_1581[31:0];
  _RAND_1582 = {1{`RANDOM}};
  stage1_regs_r_15_0_1 = _RAND_1582[31:0];
  _RAND_1583 = {1{`RANDOM}};
  stage1_regs_r_15_0_2 = _RAND_1583[31:0];
  _RAND_1584 = {1{`RANDOM}};
  stage1_regs_r_15_0_3 = _RAND_1584[31:0];
  _RAND_1585 = {1{`RANDOM}};
  stage1_regs_r_15_0_4 = _RAND_1585[31:0];
  _RAND_1586 = {1{`RANDOM}};
  stage1_regs_r_15_0_5 = _RAND_1586[31:0];
  _RAND_1587 = {1{`RANDOM}};
  stage1_regs_r_15_0_6 = _RAND_1587[31:0];
  _RAND_1588 = {1{`RANDOM}};
  stage1_regs_r_15_0_7 = _RAND_1588[31:0];
  _RAND_1589 = {1{`RANDOM}};
  stage1_regs_r_15_0_8 = _RAND_1589[31:0];
  _RAND_1590 = {1{`RANDOM}};
  stage1_regs_r_15_1_0 = _RAND_1590[31:0];
  _RAND_1591 = {1{`RANDOM}};
  stage1_regs_r_15_1_1 = _RAND_1591[31:0];
  _RAND_1592 = {1{`RANDOM}};
  stage1_regs_r_15_1_2 = _RAND_1592[31:0];
  _RAND_1593 = {1{`RANDOM}};
  stage1_regs_r_15_1_3 = _RAND_1593[31:0];
  _RAND_1594 = {1{`RANDOM}};
  stage1_regs_r_15_1_4 = _RAND_1594[31:0];
  _RAND_1595 = {1{`RANDOM}};
  stage1_regs_r_15_1_5 = _RAND_1595[31:0];
  _RAND_1596 = {1{`RANDOM}};
  stage1_regs_r_15_1_6 = _RAND_1596[31:0];
  _RAND_1597 = {1{`RANDOM}};
  stage1_regs_r_15_1_7 = _RAND_1597[31:0];
  _RAND_1598 = {1{`RANDOM}};
  stage1_regs_r_15_1_8 = _RAND_1598[31:0];
  _RAND_1599 = {1{`RANDOM}};
  stage1_regs_r_16_0_0 = _RAND_1599[31:0];
  _RAND_1600 = {1{`RANDOM}};
  stage1_regs_r_16_0_1 = _RAND_1600[31:0];
  _RAND_1601 = {1{`RANDOM}};
  stage1_regs_r_16_0_2 = _RAND_1601[31:0];
  _RAND_1602 = {1{`RANDOM}};
  stage1_regs_r_16_0_3 = _RAND_1602[31:0];
  _RAND_1603 = {1{`RANDOM}};
  stage1_regs_r_16_0_4 = _RAND_1603[31:0];
  _RAND_1604 = {1{`RANDOM}};
  stage1_regs_r_16_0_5 = _RAND_1604[31:0];
  _RAND_1605 = {1{`RANDOM}};
  stage1_regs_r_16_0_6 = _RAND_1605[31:0];
  _RAND_1606 = {1{`RANDOM}};
  stage1_regs_r_16_0_7 = _RAND_1606[31:0];
  _RAND_1607 = {1{`RANDOM}};
  stage1_regs_r_16_0_8 = _RAND_1607[31:0];
  _RAND_1608 = {1{`RANDOM}};
  stage1_regs_r_16_1_0 = _RAND_1608[31:0];
  _RAND_1609 = {1{`RANDOM}};
  stage1_regs_r_16_1_1 = _RAND_1609[31:0];
  _RAND_1610 = {1{`RANDOM}};
  stage1_regs_r_16_1_2 = _RAND_1610[31:0];
  _RAND_1611 = {1{`RANDOM}};
  stage1_regs_r_16_1_3 = _RAND_1611[31:0];
  _RAND_1612 = {1{`RANDOM}};
  stage1_regs_r_16_1_4 = _RAND_1612[31:0];
  _RAND_1613 = {1{`RANDOM}};
  stage1_regs_r_16_1_5 = _RAND_1613[31:0];
  _RAND_1614 = {1{`RANDOM}};
  stage1_regs_r_16_1_6 = _RAND_1614[31:0];
  _RAND_1615 = {1{`RANDOM}};
  stage1_regs_r_16_1_7 = _RAND_1615[31:0];
  _RAND_1616 = {1{`RANDOM}};
  stage1_regs_r_16_1_8 = _RAND_1616[31:0];
  _RAND_1617 = {1{`RANDOM}};
  stage2_regs_r_0_0_0 = _RAND_1617[31:0];
  _RAND_1618 = {1{`RANDOM}};
  stage2_regs_r_0_0_1 = _RAND_1618[31:0];
  _RAND_1619 = {1{`RANDOM}};
  stage2_regs_r_0_0_2 = _RAND_1619[31:0];
  _RAND_1620 = {1{`RANDOM}};
  stage2_regs_r_0_0_3 = _RAND_1620[31:0];
  _RAND_1621 = {1{`RANDOM}};
  stage2_regs_r_0_0_4 = _RAND_1621[31:0];
  _RAND_1622 = {1{`RANDOM}};
  stage2_regs_r_0_0_5 = _RAND_1622[31:0];
  _RAND_1623 = {1{`RANDOM}};
  stage2_regs_r_0_0_6 = _RAND_1623[31:0];
  _RAND_1624 = {1{`RANDOM}};
  stage2_regs_r_0_0_7 = _RAND_1624[31:0];
  _RAND_1625 = {1{`RANDOM}};
  stage2_regs_r_0_0_8 = _RAND_1625[31:0];
  _RAND_1626 = {1{`RANDOM}};
  stage2_regs_r_0_0_9 = _RAND_1626[31:0];
  _RAND_1627 = {1{`RANDOM}};
  stage2_regs_r_0_0_10 = _RAND_1627[31:0];
  _RAND_1628 = {1{`RANDOM}};
  stage2_regs_r_0_0_11 = _RAND_1628[31:0];
  _RAND_1629 = {1{`RANDOM}};
  stage2_regs_r_0_1_0 = _RAND_1629[31:0];
  _RAND_1630 = {1{`RANDOM}};
  stage2_regs_r_0_1_1 = _RAND_1630[31:0];
  _RAND_1631 = {1{`RANDOM}};
  stage2_regs_r_0_1_2 = _RAND_1631[31:0];
  _RAND_1632 = {1{`RANDOM}};
  stage2_regs_r_0_1_3 = _RAND_1632[31:0];
  _RAND_1633 = {1{`RANDOM}};
  stage2_regs_r_0_1_4 = _RAND_1633[31:0];
  _RAND_1634 = {1{`RANDOM}};
  stage2_regs_r_0_1_5 = _RAND_1634[31:0];
  _RAND_1635 = {1{`RANDOM}};
  stage2_regs_r_0_1_6 = _RAND_1635[31:0];
  _RAND_1636 = {1{`RANDOM}};
  stage2_regs_r_0_1_7 = _RAND_1636[31:0];
  _RAND_1637 = {1{`RANDOM}};
  stage2_regs_r_0_1_8 = _RAND_1637[31:0];
  _RAND_1638 = {1{`RANDOM}};
  stage2_regs_r_0_1_9 = _RAND_1638[31:0];
  _RAND_1639 = {1{`RANDOM}};
  stage2_regs_r_0_1_10 = _RAND_1639[31:0];
  _RAND_1640 = {1{`RANDOM}};
  stage2_regs_r_0_1_11 = _RAND_1640[31:0];
  _RAND_1641 = {1{`RANDOM}};
  stage2_regs_r_1_0_0 = _RAND_1641[31:0];
  _RAND_1642 = {1{`RANDOM}};
  stage2_regs_r_1_0_1 = _RAND_1642[31:0];
  _RAND_1643 = {1{`RANDOM}};
  stage2_regs_r_1_0_2 = _RAND_1643[31:0];
  _RAND_1644 = {1{`RANDOM}};
  stage2_regs_r_1_0_3 = _RAND_1644[31:0];
  _RAND_1645 = {1{`RANDOM}};
  stage2_regs_r_1_0_4 = _RAND_1645[31:0];
  _RAND_1646 = {1{`RANDOM}};
  stage2_regs_r_1_0_5 = _RAND_1646[31:0];
  _RAND_1647 = {1{`RANDOM}};
  stage2_regs_r_1_0_6 = _RAND_1647[31:0];
  _RAND_1648 = {1{`RANDOM}};
  stage2_regs_r_1_0_7 = _RAND_1648[31:0];
  _RAND_1649 = {1{`RANDOM}};
  stage2_regs_r_1_0_8 = _RAND_1649[31:0];
  _RAND_1650 = {1{`RANDOM}};
  stage2_regs_r_1_0_9 = _RAND_1650[31:0];
  _RAND_1651 = {1{`RANDOM}};
  stage2_regs_r_1_0_10 = _RAND_1651[31:0];
  _RAND_1652 = {1{`RANDOM}};
  stage2_regs_r_1_0_11 = _RAND_1652[31:0];
  _RAND_1653 = {1{`RANDOM}};
  stage2_regs_r_1_1_0 = _RAND_1653[31:0];
  _RAND_1654 = {1{`RANDOM}};
  stage2_regs_r_1_1_1 = _RAND_1654[31:0];
  _RAND_1655 = {1{`RANDOM}};
  stage2_regs_r_1_1_2 = _RAND_1655[31:0];
  _RAND_1656 = {1{`RANDOM}};
  stage2_regs_r_1_1_3 = _RAND_1656[31:0];
  _RAND_1657 = {1{`RANDOM}};
  stage2_regs_r_1_1_4 = _RAND_1657[31:0];
  _RAND_1658 = {1{`RANDOM}};
  stage2_regs_r_1_1_5 = _RAND_1658[31:0];
  _RAND_1659 = {1{`RANDOM}};
  stage2_regs_r_1_1_6 = _RAND_1659[31:0];
  _RAND_1660 = {1{`RANDOM}};
  stage2_regs_r_1_1_7 = _RAND_1660[31:0];
  _RAND_1661 = {1{`RANDOM}};
  stage2_regs_r_1_1_8 = _RAND_1661[31:0];
  _RAND_1662 = {1{`RANDOM}};
  stage2_regs_r_1_1_9 = _RAND_1662[31:0];
  _RAND_1663 = {1{`RANDOM}};
  stage2_regs_r_1_1_10 = _RAND_1663[31:0];
  _RAND_1664 = {1{`RANDOM}};
  stage2_regs_r_1_1_11 = _RAND_1664[31:0];
  _RAND_1665 = {1{`RANDOM}};
  stage2_regs_r_2_0_0 = _RAND_1665[31:0];
  _RAND_1666 = {1{`RANDOM}};
  stage2_regs_r_2_0_1 = _RAND_1666[31:0];
  _RAND_1667 = {1{`RANDOM}};
  stage2_regs_r_2_0_2 = _RAND_1667[31:0];
  _RAND_1668 = {1{`RANDOM}};
  stage2_regs_r_2_0_3 = _RAND_1668[31:0];
  _RAND_1669 = {1{`RANDOM}};
  stage2_regs_r_2_0_4 = _RAND_1669[31:0];
  _RAND_1670 = {1{`RANDOM}};
  stage2_regs_r_2_0_5 = _RAND_1670[31:0];
  _RAND_1671 = {1{`RANDOM}};
  stage2_regs_r_2_0_6 = _RAND_1671[31:0];
  _RAND_1672 = {1{`RANDOM}};
  stage2_regs_r_2_0_7 = _RAND_1672[31:0];
  _RAND_1673 = {1{`RANDOM}};
  stage2_regs_r_2_0_8 = _RAND_1673[31:0];
  _RAND_1674 = {1{`RANDOM}};
  stage2_regs_r_2_0_9 = _RAND_1674[31:0];
  _RAND_1675 = {1{`RANDOM}};
  stage2_regs_r_2_0_10 = _RAND_1675[31:0];
  _RAND_1676 = {1{`RANDOM}};
  stage2_regs_r_2_0_11 = _RAND_1676[31:0];
  _RAND_1677 = {1{`RANDOM}};
  stage2_regs_r_2_1_0 = _RAND_1677[31:0];
  _RAND_1678 = {1{`RANDOM}};
  stage2_regs_r_2_1_1 = _RAND_1678[31:0];
  _RAND_1679 = {1{`RANDOM}};
  stage2_regs_r_2_1_2 = _RAND_1679[31:0];
  _RAND_1680 = {1{`RANDOM}};
  stage2_regs_r_2_1_3 = _RAND_1680[31:0];
  _RAND_1681 = {1{`RANDOM}};
  stage2_regs_r_2_1_4 = _RAND_1681[31:0];
  _RAND_1682 = {1{`RANDOM}};
  stage2_regs_r_2_1_5 = _RAND_1682[31:0];
  _RAND_1683 = {1{`RANDOM}};
  stage2_regs_r_2_1_6 = _RAND_1683[31:0];
  _RAND_1684 = {1{`RANDOM}};
  stage2_regs_r_2_1_7 = _RAND_1684[31:0];
  _RAND_1685 = {1{`RANDOM}};
  stage2_regs_r_2_1_8 = _RAND_1685[31:0];
  _RAND_1686 = {1{`RANDOM}};
  stage2_regs_r_2_1_9 = _RAND_1686[31:0];
  _RAND_1687 = {1{`RANDOM}};
  stage2_regs_r_2_1_10 = _RAND_1687[31:0];
  _RAND_1688 = {1{`RANDOM}};
  stage2_regs_r_2_1_11 = _RAND_1688[31:0];
  _RAND_1689 = {1{`RANDOM}};
  stage2_regs_r_3_0_0 = _RAND_1689[31:0];
  _RAND_1690 = {1{`RANDOM}};
  stage2_regs_r_3_0_1 = _RAND_1690[31:0];
  _RAND_1691 = {1{`RANDOM}};
  stage2_regs_r_3_0_2 = _RAND_1691[31:0];
  _RAND_1692 = {1{`RANDOM}};
  stage2_regs_r_3_0_3 = _RAND_1692[31:0];
  _RAND_1693 = {1{`RANDOM}};
  stage2_regs_r_3_0_4 = _RAND_1693[31:0];
  _RAND_1694 = {1{`RANDOM}};
  stage2_regs_r_3_0_5 = _RAND_1694[31:0];
  _RAND_1695 = {1{`RANDOM}};
  stage2_regs_r_3_0_6 = _RAND_1695[31:0];
  _RAND_1696 = {1{`RANDOM}};
  stage2_regs_r_3_0_7 = _RAND_1696[31:0];
  _RAND_1697 = {1{`RANDOM}};
  stage2_regs_r_3_0_8 = _RAND_1697[31:0];
  _RAND_1698 = {1{`RANDOM}};
  stage2_regs_r_3_0_9 = _RAND_1698[31:0];
  _RAND_1699 = {1{`RANDOM}};
  stage2_regs_r_3_0_10 = _RAND_1699[31:0];
  _RAND_1700 = {1{`RANDOM}};
  stage2_regs_r_3_0_11 = _RAND_1700[31:0];
  _RAND_1701 = {1{`RANDOM}};
  stage2_regs_r_3_1_0 = _RAND_1701[31:0];
  _RAND_1702 = {1{`RANDOM}};
  stage2_regs_r_3_1_1 = _RAND_1702[31:0];
  _RAND_1703 = {1{`RANDOM}};
  stage2_regs_r_3_1_2 = _RAND_1703[31:0];
  _RAND_1704 = {1{`RANDOM}};
  stage2_regs_r_3_1_3 = _RAND_1704[31:0];
  _RAND_1705 = {1{`RANDOM}};
  stage2_regs_r_3_1_4 = _RAND_1705[31:0];
  _RAND_1706 = {1{`RANDOM}};
  stage2_regs_r_3_1_5 = _RAND_1706[31:0];
  _RAND_1707 = {1{`RANDOM}};
  stage2_regs_r_3_1_6 = _RAND_1707[31:0];
  _RAND_1708 = {1{`RANDOM}};
  stage2_regs_r_3_1_7 = _RAND_1708[31:0];
  _RAND_1709 = {1{`RANDOM}};
  stage2_regs_r_3_1_8 = _RAND_1709[31:0];
  _RAND_1710 = {1{`RANDOM}};
  stage2_regs_r_3_1_9 = _RAND_1710[31:0];
  _RAND_1711 = {1{`RANDOM}};
  stage2_regs_r_3_1_10 = _RAND_1711[31:0];
  _RAND_1712 = {1{`RANDOM}};
  stage2_regs_r_3_1_11 = _RAND_1712[31:0];
  _RAND_1713 = {1{`RANDOM}};
  stage2_regs_r_4_0_0 = _RAND_1713[31:0];
  _RAND_1714 = {1{`RANDOM}};
  stage2_regs_r_4_0_1 = _RAND_1714[31:0];
  _RAND_1715 = {1{`RANDOM}};
  stage2_regs_r_4_0_2 = _RAND_1715[31:0];
  _RAND_1716 = {1{`RANDOM}};
  stage2_regs_r_4_0_3 = _RAND_1716[31:0];
  _RAND_1717 = {1{`RANDOM}};
  stage2_regs_r_4_0_4 = _RAND_1717[31:0];
  _RAND_1718 = {1{`RANDOM}};
  stage2_regs_r_4_0_5 = _RAND_1718[31:0];
  _RAND_1719 = {1{`RANDOM}};
  stage2_regs_r_4_0_6 = _RAND_1719[31:0];
  _RAND_1720 = {1{`RANDOM}};
  stage2_regs_r_4_0_7 = _RAND_1720[31:0];
  _RAND_1721 = {1{`RANDOM}};
  stage2_regs_r_4_0_8 = _RAND_1721[31:0];
  _RAND_1722 = {1{`RANDOM}};
  stage2_regs_r_4_0_9 = _RAND_1722[31:0];
  _RAND_1723 = {1{`RANDOM}};
  stage2_regs_r_4_0_10 = _RAND_1723[31:0];
  _RAND_1724 = {1{`RANDOM}};
  stage2_regs_r_4_0_11 = _RAND_1724[31:0];
  _RAND_1725 = {1{`RANDOM}};
  stage2_regs_r_4_1_0 = _RAND_1725[31:0];
  _RAND_1726 = {1{`RANDOM}};
  stage2_regs_r_4_1_1 = _RAND_1726[31:0];
  _RAND_1727 = {1{`RANDOM}};
  stage2_regs_r_4_1_2 = _RAND_1727[31:0];
  _RAND_1728 = {1{`RANDOM}};
  stage2_regs_r_4_1_3 = _RAND_1728[31:0];
  _RAND_1729 = {1{`RANDOM}};
  stage2_regs_r_4_1_4 = _RAND_1729[31:0];
  _RAND_1730 = {1{`RANDOM}};
  stage2_regs_r_4_1_5 = _RAND_1730[31:0];
  _RAND_1731 = {1{`RANDOM}};
  stage2_regs_r_4_1_6 = _RAND_1731[31:0];
  _RAND_1732 = {1{`RANDOM}};
  stage2_regs_r_4_1_7 = _RAND_1732[31:0];
  _RAND_1733 = {1{`RANDOM}};
  stage2_regs_r_4_1_8 = _RAND_1733[31:0];
  _RAND_1734 = {1{`RANDOM}};
  stage2_regs_r_4_1_9 = _RAND_1734[31:0];
  _RAND_1735 = {1{`RANDOM}};
  stage2_regs_r_4_1_10 = _RAND_1735[31:0];
  _RAND_1736 = {1{`RANDOM}};
  stage2_regs_r_4_1_11 = _RAND_1736[31:0];
  _RAND_1737 = {1{`RANDOM}};
  stage2_regs_r_5_0_0 = _RAND_1737[31:0];
  _RAND_1738 = {1{`RANDOM}};
  stage2_regs_r_5_0_1 = _RAND_1738[31:0];
  _RAND_1739 = {1{`RANDOM}};
  stage2_regs_r_5_0_2 = _RAND_1739[31:0];
  _RAND_1740 = {1{`RANDOM}};
  stage2_regs_r_5_0_3 = _RAND_1740[31:0];
  _RAND_1741 = {1{`RANDOM}};
  stage2_regs_r_5_0_4 = _RAND_1741[31:0];
  _RAND_1742 = {1{`RANDOM}};
  stage2_regs_r_5_0_5 = _RAND_1742[31:0];
  _RAND_1743 = {1{`RANDOM}};
  stage2_regs_r_5_0_6 = _RAND_1743[31:0];
  _RAND_1744 = {1{`RANDOM}};
  stage2_regs_r_5_0_7 = _RAND_1744[31:0];
  _RAND_1745 = {1{`RANDOM}};
  stage2_regs_r_5_0_8 = _RAND_1745[31:0];
  _RAND_1746 = {1{`RANDOM}};
  stage2_regs_r_5_0_9 = _RAND_1746[31:0];
  _RAND_1747 = {1{`RANDOM}};
  stage2_regs_r_5_0_10 = _RAND_1747[31:0];
  _RAND_1748 = {1{`RANDOM}};
  stage2_regs_r_5_0_11 = _RAND_1748[31:0];
  _RAND_1749 = {1{`RANDOM}};
  stage2_regs_r_5_1_0 = _RAND_1749[31:0];
  _RAND_1750 = {1{`RANDOM}};
  stage2_regs_r_5_1_1 = _RAND_1750[31:0];
  _RAND_1751 = {1{`RANDOM}};
  stage2_regs_r_5_1_2 = _RAND_1751[31:0];
  _RAND_1752 = {1{`RANDOM}};
  stage2_regs_r_5_1_3 = _RAND_1752[31:0];
  _RAND_1753 = {1{`RANDOM}};
  stage2_regs_r_5_1_4 = _RAND_1753[31:0];
  _RAND_1754 = {1{`RANDOM}};
  stage2_regs_r_5_1_5 = _RAND_1754[31:0];
  _RAND_1755 = {1{`RANDOM}};
  stage2_regs_r_5_1_6 = _RAND_1755[31:0];
  _RAND_1756 = {1{`RANDOM}};
  stage2_regs_r_5_1_7 = _RAND_1756[31:0];
  _RAND_1757 = {1{`RANDOM}};
  stage2_regs_r_5_1_8 = _RAND_1757[31:0];
  _RAND_1758 = {1{`RANDOM}};
  stage2_regs_r_5_1_9 = _RAND_1758[31:0];
  _RAND_1759 = {1{`RANDOM}};
  stage2_regs_r_5_1_10 = _RAND_1759[31:0];
  _RAND_1760 = {1{`RANDOM}};
  stage2_regs_r_5_1_11 = _RAND_1760[31:0];
  _RAND_1761 = {1{`RANDOM}};
  stage2_regs_r_6_0_0 = _RAND_1761[31:0];
  _RAND_1762 = {1{`RANDOM}};
  stage2_regs_r_6_0_1 = _RAND_1762[31:0];
  _RAND_1763 = {1{`RANDOM}};
  stage2_regs_r_6_0_2 = _RAND_1763[31:0];
  _RAND_1764 = {1{`RANDOM}};
  stage2_regs_r_6_0_3 = _RAND_1764[31:0];
  _RAND_1765 = {1{`RANDOM}};
  stage2_regs_r_6_0_4 = _RAND_1765[31:0];
  _RAND_1766 = {1{`RANDOM}};
  stage2_regs_r_6_0_5 = _RAND_1766[31:0];
  _RAND_1767 = {1{`RANDOM}};
  stage2_regs_r_6_0_6 = _RAND_1767[31:0];
  _RAND_1768 = {1{`RANDOM}};
  stage2_regs_r_6_0_7 = _RAND_1768[31:0];
  _RAND_1769 = {1{`RANDOM}};
  stage2_regs_r_6_0_8 = _RAND_1769[31:0];
  _RAND_1770 = {1{`RANDOM}};
  stage2_regs_r_6_0_9 = _RAND_1770[31:0];
  _RAND_1771 = {1{`RANDOM}};
  stage2_regs_r_6_0_10 = _RAND_1771[31:0];
  _RAND_1772 = {1{`RANDOM}};
  stage2_regs_r_6_0_11 = _RAND_1772[31:0];
  _RAND_1773 = {1{`RANDOM}};
  stage2_regs_r_6_1_0 = _RAND_1773[31:0];
  _RAND_1774 = {1{`RANDOM}};
  stage2_regs_r_6_1_1 = _RAND_1774[31:0];
  _RAND_1775 = {1{`RANDOM}};
  stage2_regs_r_6_1_2 = _RAND_1775[31:0];
  _RAND_1776 = {1{`RANDOM}};
  stage2_regs_r_6_1_3 = _RAND_1776[31:0];
  _RAND_1777 = {1{`RANDOM}};
  stage2_regs_r_6_1_4 = _RAND_1777[31:0];
  _RAND_1778 = {1{`RANDOM}};
  stage2_regs_r_6_1_5 = _RAND_1778[31:0];
  _RAND_1779 = {1{`RANDOM}};
  stage2_regs_r_6_1_6 = _RAND_1779[31:0];
  _RAND_1780 = {1{`RANDOM}};
  stage2_regs_r_6_1_7 = _RAND_1780[31:0];
  _RAND_1781 = {1{`RANDOM}};
  stage2_regs_r_6_1_8 = _RAND_1781[31:0];
  _RAND_1782 = {1{`RANDOM}};
  stage2_regs_r_6_1_9 = _RAND_1782[31:0];
  _RAND_1783 = {1{`RANDOM}};
  stage2_regs_r_6_1_10 = _RAND_1783[31:0];
  _RAND_1784 = {1{`RANDOM}};
  stage2_regs_r_6_1_11 = _RAND_1784[31:0];
  _RAND_1785 = {1{`RANDOM}};
  stage2_regs_r_7_0_0 = _RAND_1785[31:0];
  _RAND_1786 = {1{`RANDOM}};
  stage2_regs_r_7_0_1 = _RAND_1786[31:0];
  _RAND_1787 = {1{`RANDOM}};
  stage2_regs_r_7_0_2 = _RAND_1787[31:0];
  _RAND_1788 = {1{`RANDOM}};
  stage2_regs_r_7_0_3 = _RAND_1788[31:0];
  _RAND_1789 = {1{`RANDOM}};
  stage2_regs_r_7_0_4 = _RAND_1789[31:0];
  _RAND_1790 = {1{`RANDOM}};
  stage2_regs_r_7_0_5 = _RAND_1790[31:0];
  _RAND_1791 = {1{`RANDOM}};
  stage2_regs_r_7_0_6 = _RAND_1791[31:0];
  _RAND_1792 = {1{`RANDOM}};
  stage2_regs_r_7_0_7 = _RAND_1792[31:0];
  _RAND_1793 = {1{`RANDOM}};
  stage2_regs_r_7_0_8 = _RAND_1793[31:0];
  _RAND_1794 = {1{`RANDOM}};
  stage2_regs_r_7_0_9 = _RAND_1794[31:0];
  _RAND_1795 = {1{`RANDOM}};
  stage2_regs_r_7_0_10 = _RAND_1795[31:0];
  _RAND_1796 = {1{`RANDOM}};
  stage2_regs_r_7_0_11 = _RAND_1796[31:0];
  _RAND_1797 = {1{`RANDOM}};
  stage2_regs_r_7_1_0 = _RAND_1797[31:0];
  _RAND_1798 = {1{`RANDOM}};
  stage2_regs_r_7_1_1 = _RAND_1798[31:0];
  _RAND_1799 = {1{`RANDOM}};
  stage2_regs_r_7_1_2 = _RAND_1799[31:0];
  _RAND_1800 = {1{`RANDOM}};
  stage2_regs_r_7_1_3 = _RAND_1800[31:0];
  _RAND_1801 = {1{`RANDOM}};
  stage2_regs_r_7_1_4 = _RAND_1801[31:0];
  _RAND_1802 = {1{`RANDOM}};
  stage2_regs_r_7_1_5 = _RAND_1802[31:0];
  _RAND_1803 = {1{`RANDOM}};
  stage2_regs_r_7_1_6 = _RAND_1803[31:0];
  _RAND_1804 = {1{`RANDOM}};
  stage2_regs_r_7_1_7 = _RAND_1804[31:0];
  _RAND_1805 = {1{`RANDOM}};
  stage2_regs_r_7_1_8 = _RAND_1805[31:0];
  _RAND_1806 = {1{`RANDOM}};
  stage2_regs_r_7_1_9 = _RAND_1806[31:0];
  _RAND_1807 = {1{`RANDOM}};
  stage2_regs_r_7_1_10 = _RAND_1807[31:0];
  _RAND_1808 = {1{`RANDOM}};
  stage2_regs_r_7_1_11 = _RAND_1808[31:0];
  _RAND_1809 = {1{`RANDOM}};
  stage2_regs_r_8_0_0 = _RAND_1809[31:0];
  _RAND_1810 = {1{`RANDOM}};
  stage2_regs_r_8_0_1 = _RAND_1810[31:0];
  _RAND_1811 = {1{`RANDOM}};
  stage2_regs_r_8_0_2 = _RAND_1811[31:0];
  _RAND_1812 = {1{`RANDOM}};
  stage2_regs_r_8_0_3 = _RAND_1812[31:0];
  _RAND_1813 = {1{`RANDOM}};
  stage2_regs_r_8_0_4 = _RAND_1813[31:0];
  _RAND_1814 = {1{`RANDOM}};
  stage2_regs_r_8_0_5 = _RAND_1814[31:0];
  _RAND_1815 = {1{`RANDOM}};
  stage2_regs_r_8_0_6 = _RAND_1815[31:0];
  _RAND_1816 = {1{`RANDOM}};
  stage2_regs_r_8_0_7 = _RAND_1816[31:0];
  _RAND_1817 = {1{`RANDOM}};
  stage2_regs_r_8_0_8 = _RAND_1817[31:0];
  _RAND_1818 = {1{`RANDOM}};
  stage2_regs_r_8_0_9 = _RAND_1818[31:0];
  _RAND_1819 = {1{`RANDOM}};
  stage2_regs_r_8_0_10 = _RAND_1819[31:0];
  _RAND_1820 = {1{`RANDOM}};
  stage2_regs_r_8_0_11 = _RAND_1820[31:0];
  _RAND_1821 = {1{`RANDOM}};
  stage2_regs_r_8_1_0 = _RAND_1821[31:0];
  _RAND_1822 = {1{`RANDOM}};
  stage2_regs_r_8_1_1 = _RAND_1822[31:0];
  _RAND_1823 = {1{`RANDOM}};
  stage2_regs_r_8_1_2 = _RAND_1823[31:0];
  _RAND_1824 = {1{`RANDOM}};
  stage2_regs_r_8_1_3 = _RAND_1824[31:0];
  _RAND_1825 = {1{`RANDOM}};
  stage2_regs_r_8_1_4 = _RAND_1825[31:0];
  _RAND_1826 = {1{`RANDOM}};
  stage2_regs_r_8_1_5 = _RAND_1826[31:0];
  _RAND_1827 = {1{`RANDOM}};
  stage2_regs_r_8_1_6 = _RAND_1827[31:0];
  _RAND_1828 = {1{`RANDOM}};
  stage2_regs_r_8_1_7 = _RAND_1828[31:0];
  _RAND_1829 = {1{`RANDOM}};
  stage2_regs_r_8_1_8 = _RAND_1829[31:0];
  _RAND_1830 = {1{`RANDOM}};
  stage2_regs_r_8_1_9 = _RAND_1830[31:0];
  _RAND_1831 = {1{`RANDOM}};
  stage2_regs_r_8_1_10 = _RAND_1831[31:0];
  _RAND_1832 = {1{`RANDOM}};
  stage2_regs_r_8_1_11 = _RAND_1832[31:0];
  _RAND_1833 = {1{`RANDOM}};
  stage2_regs_r_9_0_0 = _RAND_1833[31:0];
  _RAND_1834 = {1{`RANDOM}};
  stage2_regs_r_9_0_1 = _RAND_1834[31:0];
  _RAND_1835 = {1{`RANDOM}};
  stage2_regs_r_9_0_2 = _RAND_1835[31:0];
  _RAND_1836 = {1{`RANDOM}};
  stage2_regs_r_9_0_3 = _RAND_1836[31:0];
  _RAND_1837 = {1{`RANDOM}};
  stage2_regs_r_9_0_4 = _RAND_1837[31:0];
  _RAND_1838 = {1{`RANDOM}};
  stage2_regs_r_9_0_5 = _RAND_1838[31:0];
  _RAND_1839 = {1{`RANDOM}};
  stage2_regs_r_9_0_6 = _RAND_1839[31:0];
  _RAND_1840 = {1{`RANDOM}};
  stage2_regs_r_9_0_7 = _RAND_1840[31:0];
  _RAND_1841 = {1{`RANDOM}};
  stage2_regs_r_9_0_8 = _RAND_1841[31:0];
  _RAND_1842 = {1{`RANDOM}};
  stage2_regs_r_9_0_9 = _RAND_1842[31:0];
  _RAND_1843 = {1{`RANDOM}};
  stage2_regs_r_9_0_10 = _RAND_1843[31:0];
  _RAND_1844 = {1{`RANDOM}};
  stage2_regs_r_9_0_11 = _RAND_1844[31:0];
  _RAND_1845 = {1{`RANDOM}};
  stage2_regs_r_9_1_0 = _RAND_1845[31:0];
  _RAND_1846 = {1{`RANDOM}};
  stage2_regs_r_9_1_1 = _RAND_1846[31:0];
  _RAND_1847 = {1{`RANDOM}};
  stage2_regs_r_9_1_2 = _RAND_1847[31:0];
  _RAND_1848 = {1{`RANDOM}};
  stage2_regs_r_9_1_3 = _RAND_1848[31:0];
  _RAND_1849 = {1{`RANDOM}};
  stage2_regs_r_9_1_4 = _RAND_1849[31:0];
  _RAND_1850 = {1{`RANDOM}};
  stage2_regs_r_9_1_5 = _RAND_1850[31:0];
  _RAND_1851 = {1{`RANDOM}};
  stage2_regs_r_9_1_6 = _RAND_1851[31:0];
  _RAND_1852 = {1{`RANDOM}};
  stage2_regs_r_9_1_7 = _RAND_1852[31:0];
  _RAND_1853 = {1{`RANDOM}};
  stage2_regs_r_9_1_8 = _RAND_1853[31:0];
  _RAND_1854 = {1{`RANDOM}};
  stage2_regs_r_9_1_9 = _RAND_1854[31:0];
  _RAND_1855 = {1{`RANDOM}};
  stage2_regs_r_9_1_10 = _RAND_1855[31:0];
  _RAND_1856 = {1{`RANDOM}};
  stage2_regs_r_9_1_11 = _RAND_1856[31:0];
  _RAND_1857 = {1{`RANDOM}};
  stage2_regs_r_10_0_0 = _RAND_1857[31:0];
  _RAND_1858 = {1{`RANDOM}};
  stage2_regs_r_10_0_1 = _RAND_1858[31:0];
  _RAND_1859 = {1{`RANDOM}};
  stage2_regs_r_10_0_2 = _RAND_1859[31:0];
  _RAND_1860 = {1{`RANDOM}};
  stage2_regs_r_10_0_3 = _RAND_1860[31:0];
  _RAND_1861 = {1{`RANDOM}};
  stage2_regs_r_10_0_4 = _RAND_1861[31:0];
  _RAND_1862 = {1{`RANDOM}};
  stage2_regs_r_10_0_5 = _RAND_1862[31:0];
  _RAND_1863 = {1{`RANDOM}};
  stage2_regs_r_10_0_6 = _RAND_1863[31:0];
  _RAND_1864 = {1{`RANDOM}};
  stage2_regs_r_10_0_7 = _RAND_1864[31:0];
  _RAND_1865 = {1{`RANDOM}};
  stage2_regs_r_10_0_8 = _RAND_1865[31:0];
  _RAND_1866 = {1{`RANDOM}};
  stage2_regs_r_10_0_9 = _RAND_1866[31:0];
  _RAND_1867 = {1{`RANDOM}};
  stage2_regs_r_10_0_10 = _RAND_1867[31:0];
  _RAND_1868 = {1{`RANDOM}};
  stage2_regs_r_10_0_11 = _RAND_1868[31:0];
  _RAND_1869 = {1{`RANDOM}};
  stage2_regs_r_10_1_0 = _RAND_1869[31:0];
  _RAND_1870 = {1{`RANDOM}};
  stage2_regs_r_10_1_1 = _RAND_1870[31:0];
  _RAND_1871 = {1{`RANDOM}};
  stage2_regs_r_10_1_2 = _RAND_1871[31:0];
  _RAND_1872 = {1{`RANDOM}};
  stage2_regs_r_10_1_3 = _RAND_1872[31:0];
  _RAND_1873 = {1{`RANDOM}};
  stage2_regs_r_10_1_4 = _RAND_1873[31:0];
  _RAND_1874 = {1{`RANDOM}};
  stage2_regs_r_10_1_5 = _RAND_1874[31:0];
  _RAND_1875 = {1{`RANDOM}};
  stage2_regs_r_10_1_6 = _RAND_1875[31:0];
  _RAND_1876 = {1{`RANDOM}};
  stage2_regs_r_10_1_7 = _RAND_1876[31:0];
  _RAND_1877 = {1{`RANDOM}};
  stage2_regs_r_10_1_8 = _RAND_1877[31:0];
  _RAND_1878 = {1{`RANDOM}};
  stage2_regs_r_10_1_9 = _RAND_1878[31:0];
  _RAND_1879 = {1{`RANDOM}};
  stage2_regs_r_10_1_10 = _RAND_1879[31:0];
  _RAND_1880 = {1{`RANDOM}};
  stage2_regs_r_10_1_11 = _RAND_1880[31:0];
  _RAND_1881 = {1{`RANDOM}};
  stage2_regs_r_11_0_0 = _RAND_1881[31:0];
  _RAND_1882 = {1{`RANDOM}};
  stage2_regs_r_11_0_1 = _RAND_1882[31:0];
  _RAND_1883 = {1{`RANDOM}};
  stage2_regs_r_11_0_2 = _RAND_1883[31:0];
  _RAND_1884 = {1{`RANDOM}};
  stage2_regs_r_11_0_3 = _RAND_1884[31:0];
  _RAND_1885 = {1{`RANDOM}};
  stage2_regs_r_11_0_4 = _RAND_1885[31:0];
  _RAND_1886 = {1{`RANDOM}};
  stage2_regs_r_11_0_5 = _RAND_1886[31:0];
  _RAND_1887 = {1{`RANDOM}};
  stage2_regs_r_11_0_6 = _RAND_1887[31:0];
  _RAND_1888 = {1{`RANDOM}};
  stage2_regs_r_11_0_7 = _RAND_1888[31:0];
  _RAND_1889 = {1{`RANDOM}};
  stage2_regs_r_11_0_8 = _RAND_1889[31:0];
  _RAND_1890 = {1{`RANDOM}};
  stage2_regs_r_11_0_9 = _RAND_1890[31:0];
  _RAND_1891 = {1{`RANDOM}};
  stage2_regs_r_11_0_10 = _RAND_1891[31:0];
  _RAND_1892 = {1{`RANDOM}};
  stage2_regs_r_11_0_11 = _RAND_1892[31:0];
  _RAND_1893 = {1{`RANDOM}};
  stage2_regs_r_11_1_0 = _RAND_1893[31:0];
  _RAND_1894 = {1{`RANDOM}};
  stage2_regs_r_11_1_1 = _RAND_1894[31:0];
  _RAND_1895 = {1{`RANDOM}};
  stage2_regs_r_11_1_2 = _RAND_1895[31:0];
  _RAND_1896 = {1{`RANDOM}};
  stage2_regs_r_11_1_3 = _RAND_1896[31:0];
  _RAND_1897 = {1{`RANDOM}};
  stage2_regs_r_11_1_4 = _RAND_1897[31:0];
  _RAND_1898 = {1{`RANDOM}};
  stage2_regs_r_11_1_5 = _RAND_1898[31:0];
  _RAND_1899 = {1{`RANDOM}};
  stage2_regs_r_11_1_6 = _RAND_1899[31:0];
  _RAND_1900 = {1{`RANDOM}};
  stage2_regs_r_11_1_7 = _RAND_1900[31:0];
  _RAND_1901 = {1{`RANDOM}};
  stage2_regs_r_11_1_8 = _RAND_1901[31:0];
  _RAND_1902 = {1{`RANDOM}};
  stage2_regs_r_11_1_9 = _RAND_1902[31:0];
  _RAND_1903 = {1{`RANDOM}};
  stage2_regs_r_11_1_10 = _RAND_1903[31:0];
  _RAND_1904 = {1{`RANDOM}};
  stage2_regs_r_11_1_11 = _RAND_1904[31:0];
  _RAND_1905 = {1{`RANDOM}};
  stage2_regs_r_12_0_0 = _RAND_1905[31:0];
  _RAND_1906 = {1{`RANDOM}};
  stage2_regs_r_12_0_1 = _RAND_1906[31:0];
  _RAND_1907 = {1{`RANDOM}};
  stage2_regs_r_12_0_2 = _RAND_1907[31:0];
  _RAND_1908 = {1{`RANDOM}};
  stage2_regs_r_12_0_3 = _RAND_1908[31:0];
  _RAND_1909 = {1{`RANDOM}};
  stage2_regs_r_12_0_4 = _RAND_1909[31:0];
  _RAND_1910 = {1{`RANDOM}};
  stage2_regs_r_12_0_5 = _RAND_1910[31:0];
  _RAND_1911 = {1{`RANDOM}};
  stage2_regs_r_12_0_6 = _RAND_1911[31:0];
  _RAND_1912 = {1{`RANDOM}};
  stage2_regs_r_12_0_7 = _RAND_1912[31:0];
  _RAND_1913 = {1{`RANDOM}};
  stage2_regs_r_12_0_8 = _RAND_1913[31:0];
  _RAND_1914 = {1{`RANDOM}};
  stage2_regs_r_12_0_9 = _RAND_1914[31:0];
  _RAND_1915 = {1{`RANDOM}};
  stage2_regs_r_12_0_10 = _RAND_1915[31:0];
  _RAND_1916 = {1{`RANDOM}};
  stage2_regs_r_12_0_11 = _RAND_1916[31:0];
  _RAND_1917 = {1{`RANDOM}};
  stage2_regs_r_12_1_0 = _RAND_1917[31:0];
  _RAND_1918 = {1{`RANDOM}};
  stage2_regs_r_12_1_1 = _RAND_1918[31:0];
  _RAND_1919 = {1{`RANDOM}};
  stage2_regs_r_12_1_2 = _RAND_1919[31:0];
  _RAND_1920 = {1{`RANDOM}};
  stage2_regs_r_12_1_3 = _RAND_1920[31:0];
  _RAND_1921 = {1{`RANDOM}};
  stage2_regs_r_12_1_4 = _RAND_1921[31:0];
  _RAND_1922 = {1{`RANDOM}};
  stage2_regs_r_12_1_5 = _RAND_1922[31:0];
  _RAND_1923 = {1{`RANDOM}};
  stage2_regs_r_12_1_6 = _RAND_1923[31:0];
  _RAND_1924 = {1{`RANDOM}};
  stage2_regs_r_12_1_7 = _RAND_1924[31:0];
  _RAND_1925 = {1{`RANDOM}};
  stage2_regs_r_12_1_8 = _RAND_1925[31:0];
  _RAND_1926 = {1{`RANDOM}};
  stage2_regs_r_12_1_9 = _RAND_1926[31:0];
  _RAND_1927 = {1{`RANDOM}};
  stage2_regs_r_12_1_10 = _RAND_1927[31:0];
  _RAND_1928 = {1{`RANDOM}};
  stage2_regs_r_12_1_11 = _RAND_1928[31:0];
  _RAND_1929 = {1{`RANDOM}};
  stage2_regs_r_13_0_0 = _RAND_1929[31:0];
  _RAND_1930 = {1{`RANDOM}};
  stage2_regs_r_13_0_1 = _RAND_1930[31:0];
  _RAND_1931 = {1{`RANDOM}};
  stage2_regs_r_13_0_2 = _RAND_1931[31:0];
  _RAND_1932 = {1{`RANDOM}};
  stage2_regs_r_13_0_3 = _RAND_1932[31:0];
  _RAND_1933 = {1{`RANDOM}};
  stage2_regs_r_13_0_4 = _RAND_1933[31:0];
  _RAND_1934 = {1{`RANDOM}};
  stage2_regs_r_13_0_5 = _RAND_1934[31:0];
  _RAND_1935 = {1{`RANDOM}};
  stage2_regs_r_13_0_6 = _RAND_1935[31:0];
  _RAND_1936 = {1{`RANDOM}};
  stage2_regs_r_13_0_7 = _RAND_1936[31:0];
  _RAND_1937 = {1{`RANDOM}};
  stage2_regs_r_13_0_8 = _RAND_1937[31:0];
  _RAND_1938 = {1{`RANDOM}};
  stage2_regs_r_13_0_9 = _RAND_1938[31:0];
  _RAND_1939 = {1{`RANDOM}};
  stage2_regs_r_13_0_10 = _RAND_1939[31:0];
  _RAND_1940 = {1{`RANDOM}};
  stage2_regs_r_13_0_11 = _RAND_1940[31:0];
  _RAND_1941 = {1{`RANDOM}};
  stage2_regs_r_13_1_0 = _RAND_1941[31:0];
  _RAND_1942 = {1{`RANDOM}};
  stage2_regs_r_13_1_1 = _RAND_1942[31:0];
  _RAND_1943 = {1{`RANDOM}};
  stage2_regs_r_13_1_2 = _RAND_1943[31:0];
  _RAND_1944 = {1{`RANDOM}};
  stage2_regs_r_13_1_3 = _RAND_1944[31:0];
  _RAND_1945 = {1{`RANDOM}};
  stage2_regs_r_13_1_4 = _RAND_1945[31:0];
  _RAND_1946 = {1{`RANDOM}};
  stage2_regs_r_13_1_5 = _RAND_1946[31:0];
  _RAND_1947 = {1{`RANDOM}};
  stage2_regs_r_13_1_6 = _RAND_1947[31:0];
  _RAND_1948 = {1{`RANDOM}};
  stage2_regs_r_13_1_7 = _RAND_1948[31:0];
  _RAND_1949 = {1{`RANDOM}};
  stage2_regs_r_13_1_8 = _RAND_1949[31:0];
  _RAND_1950 = {1{`RANDOM}};
  stage2_regs_r_13_1_9 = _RAND_1950[31:0];
  _RAND_1951 = {1{`RANDOM}};
  stage2_regs_r_13_1_10 = _RAND_1951[31:0];
  _RAND_1952 = {1{`RANDOM}};
  stage2_regs_r_13_1_11 = _RAND_1952[31:0];
  _RAND_1953 = {1{`RANDOM}};
  stage2_regs_r_14_0_0 = _RAND_1953[31:0];
  _RAND_1954 = {1{`RANDOM}};
  stage2_regs_r_14_0_1 = _RAND_1954[31:0];
  _RAND_1955 = {1{`RANDOM}};
  stage2_regs_r_14_0_2 = _RAND_1955[31:0];
  _RAND_1956 = {1{`RANDOM}};
  stage2_regs_r_14_0_3 = _RAND_1956[31:0];
  _RAND_1957 = {1{`RANDOM}};
  stage2_regs_r_14_0_4 = _RAND_1957[31:0];
  _RAND_1958 = {1{`RANDOM}};
  stage2_regs_r_14_0_5 = _RAND_1958[31:0];
  _RAND_1959 = {1{`RANDOM}};
  stage2_regs_r_14_0_6 = _RAND_1959[31:0];
  _RAND_1960 = {1{`RANDOM}};
  stage2_regs_r_14_0_7 = _RAND_1960[31:0];
  _RAND_1961 = {1{`RANDOM}};
  stage2_regs_r_14_0_8 = _RAND_1961[31:0];
  _RAND_1962 = {1{`RANDOM}};
  stage2_regs_r_14_0_9 = _RAND_1962[31:0];
  _RAND_1963 = {1{`RANDOM}};
  stage2_regs_r_14_0_10 = _RAND_1963[31:0];
  _RAND_1964 = {1{`RANDOM}};
  stage2_regs_r_14_0_11 = _RAND_1964[31:0];
  _RAND_1965 = {1{`RANDOM}};
  stage2_regs_r_14_1_0 = _RAND_1965[31:0];
  _RAND_1966 = {1{`RANDOM}};
  stage2_regs_r_14_1_1 = _RAND_1966[31:0];
  _RAND_1967 = {1{`RANDOM}};
  stage2_regs_r_14_1_2 = _RAND_1967[31:0];
  _RAND_1968 = {1{`RANDOM}};
  stage2_regs_r_14_1_3 = _RAND_1968[31:0];
  _RAND_1969 = {1{`RANDOM}};
  stage2_regs_r_14_1_4 = _RAND_1969[31:0];
  _RAND_1970 = {1{`RANDOM}};
  stage2_regs_r_14_1_5 = _RAND_1970[31:0];
  _RAND_1971 = {1{`RANDOM}};
  stage2_regs_r_14_1_6 = _RAND_1971[31:0];
  _RAND_1972 = {1{`RANDOM}};
  stage2_regs_r_14_1_7 = _RAND_1972[31:0];
  _RAND_1973 = {1{`RANDOM}};
  stage2_regs_r_14_1_8 = _RAND_1973[31:0];
  _RAND_1974 = {1{`RANDOM}};
  stage2_regs_r_14_1_9 = _RAND_1974[31:0];
  _RAND_1975 = {1{`RANDOM}};
  stage2_regs_r_14_1_10 = _RAND_1975[31:0];
  _RAND_1976 = {1{`RANDOM}};
  stage2_regs_r_14_1_11 = _RAND_1976[31:0];
  _RAND_1977 = {1{`RANDOM}};
  stage2_regs_r_15_0_0 = _RAND_1977[31:0];
  _RAND_1978 = {1{`RANDOM}};
  stage2_regs_r_15_0_1 = _RAND_1978[31:0];
  _RAND_1979 = {1{`RANDOM}};
  stage2_regs_r_15_0_2 = _RAND_1979[31:0];
  _RAND_1980 = {1{`RANDOM}};
  stage2_regs_r_15_0_3 = _RAND_1980[31:0];
  _RAND_1981 = {1{`RANDOM}};
  stage2_regs_r_15_0_4 = _RAND_1981[31:0];
  _RAND_1982 = {1{`RANDOM}};
  stage2_regs_r_15_0_5 = _RAND_1982[31:0];
  _RAND_1983 = {1{`RANDOM}};
  stage2_regs_r_15_0_6 = _RAND_1983[31:0];
  _RAND_1984 = {1{`RANDOM}};
  stage2_regs_r_15_0_7 = _RAND_1984[31:0];
  _RAND_1985 = {1{`RANDOM}};
  stage2_regs_r_15_0_8 = _RAND_1985[31:0];
  _RAND_1986 = {1{`RANDOM}};
  stage2_regs_r_15_0_9 = _RAND_1986[31:0];
  _RAND_1987 = {1{`RANDOM}};
  stage2_regs_r_15_0_10 = _RAND_1987[31:0];
  _RAND_1988 = {1{`RANDOM}};
  stage2_regs_r_15_0_11 = _RAND_1988[31:0];
  _RAND_1989 = {1{`RANDOM}};
  stage2_regs_r_15_1_0 = _RAND_1989[31:0];
  _RAND_1990 = {1{`RANDOM}};
  stage2_regs_r_15_1_1 = _RAND_1990[31:0];
  _RAND_1991 = {1{`RANDOM}};
  stage2_regs_r_15_1_2 = _RAND_1991[31:0];
  _RAND_1992 = {1{`RANDOM}};
  stage2_regs_r_15_1_3 = _RAND_1992[31:0];
  _RAND_1993 = {1{`RANDOM}};
  stage2_regs_r_15_1_4 = _RAND_1993[31:0];
  _RAND_1994 = {1{`RANDOM}};
  stage2_regs_r_15_1_5 = _RAND_1994[31:0];
  _RAND_1995 = {1{`RANDOM}};
  stage2_regs_r_15_1_6 = _RAND_1995[31:0];
  _RAND_1996 = {1{`RANDOM}};
  stage2_regs_r_15_1_7 = _RAND_1996[31:0];
  _RAND_1997 = {1{`RANDOM}};
  stage2_regs_r_15_1_8 = _RAND_1997[31:0];
  _RAND_1998 = {1{`RANDOM}};
  stage2_regs_r_15_1_9 = _RAND_1998[31:0];
  _RAND_1999 = {1{`RANDOM}};
  stage2_regs_r_15_1_10 = _RAND_1999[31:0];
  _RAND_2000 = {1{`RANDOM}};
  stage2_regs_r_15_1_11 = _RAND_2000[31:0];
  _RAND_2001 = {1{`RANDOM}};
  stage2_regs_r_16_0_0 = _RAND_2001[31:0];
  _RAND_2002 = {1{`RANDOM}};
  stage2_regs_r_16_0_1 = _RAND_2002[31:0];
  _RAND_2003 = {1{`RANDOM}};
  stage2_regs_r_16_0_2 = _RAND_2003[31:0];
  _RAND_2004 = {1{`RANDOM}};
  stage2_regs_r_16_0_3 = _RAND_2004[31:0];
  _RAND_2005 = {1{`RANDOM}};
  stage2_regs_r_16_0_4 = _RAND_2005[31:0];
  _RAND_2006 = {1{`RANDOM}};
  stage2_regs_r_16_0_5 = _RAND_2006[31:0];
  _RAND_2007 = {1{`RANDOM}};
  stage2_regs_r_16_0_6 = _RAND_2007[31:0];
  _RAND_2008 = {1{`RANDOM}};
  stage2_regs_r_16_0_7 = _RAND_2008[31:0];
  _RAND_2009 = {1{`RANDOM}};
  stage2_regs_r_16_0_8 = _RAND_2009[31:0];
  _RAND_2010 = {1{`RANDOM}};
  stage2_regs_r_16_0_9 = _RAND_2010[31:0];
  _RAND_2011 = {1{`RANDOM}};
  stage2_regs_r_16_0_10 = _RAND_2011[31:0];
  _RAND_2012 = {1{`RANDOM}};
  stage2_regs_r_16_0_11 = _RAND_2012[31:0];
  _RAND_2013 = {1{`RANDOM}};
  stage2_regs_r_16_1_0 = _RAND_2013[31:0];
  _RAND_2014 = {1{`RANDOM}};
  stage2_regs_r_16_1_1 = _RAND_2014[31:0];
  _RAND_2015 = {1{`RANDOM}};
  stage2_regs_r_16_1_2 = _RAND_2015[31:0];
  _RAND_2016 = {1{`RANDOM}};
  stage2_regs_r_16_1_3 = _RAND_2016[31:0];
  _RAND_2017 = {1{`RANDOM}};
  stage2_regs_r_16_1_4 = _RAND_2017[31:0];
  _RAND_2018 = {1{`RANDOM}};
  stage2_regs_r_16_1_5 = _RAND_2018[31:0];
  _RAND_2019 = {1{`RANDOM}};
  stage2_regs_r_16_1_6 = _RAND_2019[31:0];
  _RAND_2020 = {1{`RANDOM}};
  stage2_regs_r_16_1_7 = _RAND_2020[31:0];
  _RAND_2021 = {1{`RANDOM}};
  stage2_regs_r_16_1_8 = _RAND_2021[31:0];
  _RAND_2022 = {1{`RANDOM}};
  stage2_regs_r_16_1_9 = _RAND_2022[31:0];
  _RAND_2023 = {1{`RANDOM}};
  stage2_regs_r_16_1_10 = _RAND_2023[31:0];
  _RAND_2024 = {1{`RANDOM}};
  stage2_regs_r_16_1_11 = _RAND_2024[31:0];
  _RAND_2025 = {1{`RANDOM}};
  stage3_regs_r_0_1_0 = _RAND_2025[31:0];
  _RAND_2026 = {1{`RANDOM}};
  stage3_regs_r_0_1_1 = _RAND_2026[31:0];
  _RAND_2027 = {1{`RANDOM}};
  stage3_regs_r_0_1_2 = _RAND_2027[31:0];
  _RAND_2028 = {1{`RANDOM}};
  stage3_regs_r_0_1_3 = _RAND_2028[31:0];
  _RAND_2029 = {1{`RANDOM}};
  stage3_regs_r_0_1_4 = _RAND_2029[31:0];
  _RAND_2030 = {1{`RANDOM}};
  stage3_regs_r_0_1_5 = _RAND_2030[31:0];
  _RAND_2031 = {1{`RANDOM}};
  stage3_regs_r_0_1_6 = _RAND_2031[31:0];
  _RAND_2032 = {1{`RANDOM}};
  stage3_regs_r_0_1_7 = _RAND_2032[31:0];
  _RAND_2033 = {1{`RANDOM}};
  stage3_regs_r_0_1_8 = _RAND_2033[31:0];
  _RAND_2034 = {1{`RANDOM}};
  stage3_regs_r_1_1_0 = _RAND_2034[31:0];
  _RAND_2035 = {1{`RANDOM}};
  stage3_regs_r_1_1_1 = _RAND_2035[31:0];
  _RAND_2036 = {1{`RANDOM}};
  stage3_regs_r_1_1_2 = _RAND_2036[31:0];
  _RAND_2037 = {1{`RANDOM}};
  stage3_regs_r_1_1_3 = _RAND_2037[31:0];
  _RAND_2038 = {1{`RANDOM}};
  stage3_regs_r_1_1_4 = _RAND_2038[31:0];
  _RAND_2039 = {1{`RANDOM}};
  stage3_regs_r_1_1_5 = _RAND_2039[31:0];
  _RAND_2040 = {1{`RANDOM}};
  stage3_regs_r_1_1_6 = _RAND_2040[31:0];
  _RAND_2041 = {1{`RANDOM}};
  stage3_regs_r_1_1_7 = _RAND_2041[31:0];
  _RAND_2042 = {1{`RANDOM}};
  stage3_regs_r_1_1_8 = _RAND_2042[31:0];
  _RAND_2043 = {1{`RANDOM}};
  stage3_regs_r_2_1_0 = _RAND_2043[31:0];
  _RAND_2044 = {1{`RANDOM}};
  stage3_regs_r_2_1_1 = _RAND_2044[31:0];
  _RAND_2045 = {1{`RANDOM}};
  stage3_regs_r_2_1_2 = _RAND_2045[31:0];
  _RAND_2046 = {1{`RANDOM}};
  stage3_regs_r_2_1_3 = _RAND_2046[31:0];
  _RAND_2047 = {1{`RANDOM}};
  stage3_regs_r_2_1_4 = _RAND_2047[31:0];
  _RAND_2048 = {1{`RANDOM}};
  stage3_regs_r_2_1_5 = _RAND_2048[31:0];
  _RAND_2049 = {1{`RANDOM}};
  stage3_regs_r_2_1_6 = _RAND_2049[31:0];
  _RAND_2050 = {1{`RANDOM}};
  stage3_regs_r_2_1_7 = _RAND_2050[31:0];
  _RAND_2051 = {1{`RANDOM}};
  stage3_regs_r_2_1_8 = _RAND_2051[31:0];
  _RAND_2052 = {1{`RANDOM}};
  stage3_regs_r_3_1_0 = _RAND_2052[31:0];
  _RAND_2053 = {1{`RANDOM}};
  stage3_regs_r_3_1_1 = _RAND_2053[31:0];
  _RAND_2054 = {1{`RANDOM}};
  stage3_regs_r_3_1_2 = _RAND_2054[31:0];
  _RAND_2055 = {1{`RANDOM}};
  stage3_regs_r_3_1_3 = _RAND_2055[31:0];
  _RAND_2056 = {1{`RANDOM}};
  stage3_regs_r_3_1_4 = _RAND_2056[31:0];
  _RAND_2057 = {1{`RANDOM}};
  stage3_regs_r_3_1_5 = _RAND_2057[31:0];
  _RAND_2058 = {1{`RANDOM}};
  stage3_regs_r_3_1_6 = _RAND_2058[31:0];
  _RAND_2059 = {1{`RANDOM}};
  stage3_regs_r_3_1_7 = _RAND_2059[31:0];
  _RAND_2060 = {1{`RANDOM}};
  stage3_regs_r_3_1_8 = _RAND_2060[31:0];
  _RAND_2061 = {1{`RANDOM}};
  stage3_regs_r_4_1_0 = _RAND_2061[31:0];
  _RAND_2062 = {1{`RANDOM}};
  stage3_regs_r_4_1_1 = _RAND_2062[31:0];
  _RAND_2063 = {1{`RANDOM}};
  stage3_regs_r_4_1_2 = _RAND_2063[31:0];
  _RAND_2064 = {1{`RANDOM}};
  stage3_regs_r_4_1_3 = _RAND_2064[31:0];
  _RAND_2065 = {1{`RANDOM}};
  stage3_regs_r_4_1_4 = _RAND_2065[31:0];
  _RAND_2066 = {1{`RANDOM}};
  stage3_regs_r_4_1_5 = _RAND_2066[31:0];
  _RAND_2067 = {1{`RANDOM}};
  stage3_regs_r_4_1_6 = _RAND_2067[31:0];
  _RAND_2068 = {1{`RANDOM}};
  stage3_regs_r_4_1_7 = _RAND_2068[31:0];
  _RAND_2069 = {1{`RANDOM}};
  stage3_regs_r_4_1_8 = _RAND_2069[31:0];
  _RAND_2070 = {1{`RANDOM}};
  stage3_regs_r_5_1_0 = _RAND_2070[31:0];
  _RAND_2071 = {1{`RANDOM}};
  stage3_regs_r_5_1_1 = _RAND_2071[31:0];
  _RAND_2072 = {1{`RANDOM}};
  stage3_regs_r_5_1_2 = _RAND_2072[31:0];
  _RAND_2073 = {1{`RANDOM}};
  stage3_regs_r_5_1_3 = _RAND_2073[31:0];
  _RAND_2074 = {1{`RANDOM}};
  stage3_regs_r_5_1_4 = _RAND_2074[31:0];
  _RAND_2075 = {1{`RANDOM}};
  stage3_regs_r_5_1_5 = _RAND_2075[31:0];
  _RAND_2076 = {1{`RANDOM}};
  stage3_regs_r_5_1_6 = _RAND_2076[31:0];
  _RAND_2077 = {1{`RANDOM}};
  stage3_regs_r_5_1_7 = _RAND_2077[31:0];
  _RAND_2078 = {1{`RANDOM}};
  stage3_regs_r_5_1_8 = _RAND_2078[31:0];
  _RAND_2079 = {1{`RANDOM}};
  stage3_regs_r_6_1_0 = _RAND_2079[31:0];
  _RAND_2080 = {1{`RANDOM}};
  stage3_regs_r_6_1_1 = _RAND_2080[31:0];
  _RAND_2081 = {1{`RANDOM}};
  stage3_regs_r_6_1_2 = _RAND_2081[31:0];
  _RAND_2082 = {1{`RANDOM}};
  stage3_regs_r_6_1_3 = _RAND_2082[31:0];
  _RAND_2083 = {1{`RANDOM}};
  stage3_regs_r_6_1_4 = _RAND_2083[31:0];
  _RAND_2084 = {1{`RANDOM}};
  stage3_regs_r_6_1_5 = _RAND_2084[31:0];
  _RAND_2085 = {1{`RANDOM}};
  stage3_regs_r_6_1_6 = _RAND_2085[31:0];
  _RAND_2086 = {1{`RANDOM}};
  stage3_regs_r_6_1_7 = _RAND_2086[31:0];
  _RAND_2087 = {1{`RANDOM}};
  stage3_regs_r_6_1_8 = _RAND_2087[31:0];
  _RAND_2088 = {1{`RANDOM}};
  stage3_regs_r_7_1_0 = _RAND_2088[31:0];
  _RAND_2089 = {1{`RANDOM}};
  stage3_regs_r_7_1_1 = _RAND_2089[31:0];
  _RAND_2090 = {1{`RANDOM}};
  stage3_regs_r_7_1_2 = _RAND_2090[31:0];
  _RAND_2091 = {1{`RANDOM}};
  stage3_regs_r_7_1_3 = _RAND_2091[31:0];
  _RAND_2092 = {1{`RANDOM}};
  stage3_regs_r_7_1_4 = _RAND_2092[31:0];
  _RAND_2093 = {1{`RANDOM}};
  stage3_regs_r_7_1_5 = _RAND_2093[31:0];
  _RAND_2094 = {1{`RANDOM}};
  stage3_regs_r_7_1_6 = _RAND_2094[31:0];
  _RAND_2095 = {1{`RANDOM}};
  stage3_regs_r_7_1_7 = _RAND_2095[31:0];
  _RAND_2096 = {1{`RANDOM}};
  stage3_regs_r_7_1_8 = _RAND_2096[31:0];
  _RAND_2097 = {1{`RANDOM}};
  stage3_regs_r_8_1_0 = _RAND_2097[31:0];
  _RAND_2098 = {1{`RANDOM}};
  stage3_regs_r_8_1_1 = _RAND_2098[31:0];
  _RAND_2099 = {1{`RANDOM}};
  stage3_regs_r_8_1_2 = _RAND_2099[31:0];
  _RAND_2100 = {1{`RANDOM}};
  stage3_regs_r_8_1_3 = _RAND_2100[31:0];
  _RAND_2101 = {1{`RANDOM}};
  stage3_regs_r_8_1_4 = _RAND_2101[31:0];
  _RAND_2102 = {1{`RANDOM}};
  stage3_regs_r_8_1_5 = _RAND_2102[31:0];
  _RAND_2103 = {1{`RANDOM}};
  stage3_regs_r_8_1_6 = _RAND_2103[31:0];
  _RAND_2104 = {1{`RANDOM}};
  stage3_regs_r_8_1_7 = _RAND_2104[31:0];
  _RAND_2105 = {1{`RANDOM}};
  stage3_regs_r_8_1_8 = _RAND_2105[31:0];
  _RAND_2106 = {1{`RANDOM}};
  stage3_regs_r_9_1_0 = _RAND_2106[31:0];
  _RAND_2107 = {1{`RANDOM}};
  stage3_regs_r_9_1_1 = _RAND_2107[31:0];
  _RAND_2108 = {1{`RANDOM}};
  stage3_regs_r_9_1_2 = _RAND_2108[31:0];
  _RAND_2109 = {1{`RANDOM}};
  stage3_regs_r_9_1_3 = _RAND_2109[31:0];
  _RAND_2110 = {1{`RANDOM}};
  stage3_regs_r_9_1_4 = _RAND_2110[31:0];
  _RAND_2111 = {1{`RANDOM}};
  stage3_regs_r_9_1_5 = _RAND_2111[31:0];
  _RAND_2112 = {1{`RANDOM}};
  stage3_regs_r_9_1_6 = _RAND_2112[31:0];
  _RAND_2113 = {1{`RANDOM}};
  stage3_regs_r_9_1_7 = _RAND_2113[31:0];
  _RAND_2114 = {1{`RANDOM}};
  stage3_regs_r_9_1_8 = _RAND_2114[31:0];
  _RAND_2115 = {1{`RANDOM}};
  stage3_regs_r_10_1_0 = _RAND_2115[31:0];
  _RAND_2116 = {1{`RANDOM}};
  stage3_regs_r_10_1_1 = _RAND_2116[31:0];
  _RAND_2117 = {1{`RANDOM}};
  stage3_regs_r_10_1_2 = _RAND_2117[31:0];
  _RAND_2118 = {1{`RANDOM}};
  stage3_regs_r_10_1_3 = _RAND_2118[31:0];
  _RAND_2119 = {1{`RANDOM}};
  stage3_regs_r_10_1_4 = _RAND_2119[31:0];
  _RAND_2120 = {1{`RANDOM}};
  stage3_regs_r_10_1_5 = _RAND_2120[31:0];
  _RAND_2121 = {1{`RANDOM}};
  stage3_regs_r_10_1_6 = _RAND_2121[31:0];
  _RAND_2122 = {1{`RANDOM}};
  stage3_regs_r_10_1_7 = _RAND_2122[31:0];
  _RAND_2123 = {1{`RANDOM}};
  stage3_regs_r_10_1_8 = _RAND_2123[31:0];
  _RAND_2124 = {1{`RANDOM}};
  stage3_regs_r_11_1_0 = _RAND_2124[31:0];
  _RAND_2125 = {1{`RANDOM}};
  stage3_regs_r_11_1_1 = _RAND_2125[31:0];
  _RAND_2126 = {1{`RANDOM}};
  stage3_regs_r_11_1_2 = _RAND_2126[31:0];
  _RAND_2127 = {1{`RANDOM}};
  stage3_regs_r_11_1_3 = _RAND_2127[31:0];
  _RAND_2128 = {1{`RANDOM}};
  stage3_regs_r_11_1_4 = _RAND_2128[31:0];
  _RAND_2129 = {1{`RANDOM}};
  stage3_regs_r_11_1_5 = _RAND_2129[31:0];
  _RAND_2130 = {1{`RANDOM}};
  stage3_regs_r_11_1_6 = _RAND_2130[31:0];
  _RAND_2131 = {1{`RANDOM}};
  stage3_regs_r_11_1_7 = _RAND_2131[31:0];
  _RAND_2132 = {1{`RANDOM}};
  stage3_regs_r_11_1_8 = _RAND_2132[31:0];
  _RAND_2133 = {1{`RANDOM}};
  stage3_regs_r_12_1_0 = _RAND_2133[31:0];
  _RAND_2134 = {1{`RANDOM}};
  stage3_regs_r_12_1_1 = _RAND_2134[31:0];
  _RAND_2135 = {1{`RANDOM}};
  stage3_regs_r_12_1_2 = _RAND_2135[31:0];
  _RAND_2136 = {1{`RANDOM}};
  stage3_regs_r_12_1_3 = _RAND_2136[31:0];
  _RAND_2137 = {1{`RANDOM}};
  stage3_regs_r_12_1_4 = _RAND_2137[31:0];
  _RAND_2138 = {1{`RANDOM}};
  stage3_regs_r_12_1_5 = _RAND_2138[31:0];
  _RAND_2139 = {1{`RANDOM}};
  stage3_regs_r_12_1_6 = _RAND_2139[31:0];
  _RAND_2140 = {1{`RANDOM}};
  stage3_regs_r_12_1_7 = _RAND_2140[31:0];
  _RAND_2141 = {1{`RANDOM}};
  stage3_regs_r_12_1_8 = _RAND_2141[31:0];
  _RAND_2142 = {1{`RANDOM}};
  stage3_regs_r_13_1_0 = _RAND_2142[31:0];
  _RAND_2143 = {1{`RANDOM}};
  stage3_regs_r_13_1_1 = _RAND_2143[31:0];
  _RAND_2144 = {1{`RANDOM}};
  stage3_regs_r_13_1_2 = _RAND_2144[31:0];
  _RAND_2145 = {1{`RANDOM}};
  stage3_regs_r_13_1_3 = _RAND_2145[31:0];
  _RAND_2146 = {1{`RANDOM}};
  stage3_regs_r_13_1_4 = _RAND_2146[31:0];
  _RAND_2147 = {1{`RANDOM}};
  stage3_regs_r_13_1_5 = _RAND_2147[31:0];
  _RAND_2148 = {1{`RANDOM}};
  stage3_regs_r_13_1_6 = _RAND_2148[31:0];
  _RAND_2149 = {1{`RANDOM}};
  stage3_regs_r_13_1_7 = _RAND_2149[31:0];
  _RAND_2150 = {1{`RANDOM}};
  stage3_regs_r_13_1_8 = _RAND_2150[31:0];
  _RAND_2151 = {1{`RANDOM}};
  stage3_regs_r_14_1_0 = _RAND_2151[31:0];
  _RAND_2152 = {1{`RANDOM}};
  stage3_regs_r_14_1_1 = _RAND_2152[31:0];
  _RAND_2153 = {1{`RANDOM}};
  stage3_regs_r_14_1_2 = _RAND_2153[31:0];
  _RAND_2154 = {1{`RANDOM}};
  stage3_regs_r_14_1_3 = _RAND_2154[31:0];
  _RAND_2155 = {1{`RANDOM}};
  stage3_regs_r_14_1_4 = _RAND_2155[31:0];
  _RAND_2156 = {1{`RANDOM}};
  stage3_regs_r_14_1_5 = _RAND_2156[31:0];
  _RAND_2157 = {1{`RANDOM}};
  stage3_regs_r_14_1_6 = _RAND_2157[31:0];
  _RAND_2158 = {1{`RANDOM}};
  stage3_regs_r_14_1_7 = _RAND_2158[31:0];
  _RAND_2159 = {1{`RANDOM}};
  stage3_regs_r_14_1_8 = _RAND_2159[31:0];
  _RAND_2160 = {1{`RANDOM}};
  stage3_regs_r_15_1_0 = _RAND_2160[31:0];
  _RAND_2161 = {1{`RANDOM}};
  stage3_regs_r_15_1_1 = _RAND_2161[31:0];
  _RAND_2162 = {1{`RANDOM}};
  stage3_regs_r_15_1_2 = _RAND_2162[31:0];
  _RAND_2163 = {1{`RANDOM}};
  stage3_regs_r_15_1_3 = _RAND_2163[31:0];
  _RAND_2164 = {1{`RANDOM}};
  stage3_regs_r_15_1_4 = _RAND_2164[31:0];
  _RAND_2165 = {1{`RANDOM}};
  stage3_regs_r_15_1_5 = _RAND_2165[31:0];
  _RAND_2166 = {1{`RANDOM}};
  stage3_regs_r_15_1_6 = _RAND_2166[31:0];
  _RAND_2167 = {1{`RANDOM}};
  stage3_regs_r_15_1_7 = _RAND_2167[31:0];
  _RAND_2168 = {1{`RANDOM}};
  stage3_regs_r_15_1_8 = _RAND_2168[31:0];
  _RAND_2169 = {1{`RANDOM}};
  stage3_regs_r_16_1_0 = _RAND_2169[31:0];
  _RAND_2170 = {1{`RANDOM}};
  stage3_regs_r_16_1_1 = _RAND_2170[31:0];
  _RAND_2171 = {1{`RANDOM}};
  stage3_regs_r_16_1_2 = _RAND_2171[31:0];
  _RAND_2172 = {1{`RANDOM}};
  stage3_regs_r_16_1_3 = _RAND_2172[31:0];
  _RAND_2173 = {1{`RANDOM}};
  stage3_regs_r_16_1_4 = _RAND_2173[31:0];
  _RAND_2174 = {1{`RANDOM}};
  stage3_regs_r_16_1_5 = _RAND_2174[31:0];
  _RAND_2175 = {1{`RANDOM}};
  stage3_regs_r_16_1_6 = _RAND_2175[31:0];
  _RAND_2176 = {1{`RANDOM}};
  stage3_regs_r_16_1_7 = _RAND_2176[31:0];
  _RAND_2177 = {1{`RANDOM}};
  stage3_regs_r_16_1_8 = _RAND_2177[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FP_divider_newfpu(
  input         clock,
  input         reset,
  input         io_in_en,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
`endif // RANDOMIZE_REG_INIT
  wire  FP_reciprocal_newfpu_clock; // @[FloatingPointDesigns.scala 2279:28]
  wire  FP_reciprocal_newfpu_reset; // @[FloatingPointDesigns.scala 2279:28]
  wire  FP_reciprocal_newfpu_io_in_en; // @[FloatingPointDesigns.scala 2279:28]
  wire [31:0] FP_reciprocal_newfpu_io_in_a; // @[FloatingPointDesigns.scala 2279:28]
  wire [31:0] FP_reciprocal_newfpu_io_out_s; // @[FloatingPointDesigns.scala 2279:28]
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 2282:28]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 2282:28]
  wire  FP_multiplier_10ccs_io_in_en; // @[FloatingPointDesigns.scala 2282:28]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 2282:28]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 2282:28]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2282:28]
  reg [31:0] regs_0; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_2; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_3; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_4; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_5; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_6; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_7; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_8; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_9; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_10; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_11; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_12; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_13; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_14; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_15; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_16; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_17; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_18; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_19; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_20; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_21; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_22; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_23; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_24; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_25; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_26; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_27; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_28; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_29; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_30; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_31; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_32; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_33; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_34; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_35; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_36; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_37; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_38; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_39; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_40; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_41; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_42; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_43; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_44; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_45; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_46; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_47; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_48; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_49; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_50; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_51; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_52; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_53; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_54; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_55; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_56; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_57; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_58; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_59; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_60; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_61; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_62; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_63; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_64; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_65; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_66; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_67; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_68; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_69; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_70; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_71; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_72; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_73; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_74; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_75; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_76; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_77; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_78; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_79; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_80; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_81; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_82; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_83; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_84; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_85; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_86; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_87; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_88; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_89; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_90; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_91; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_92; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_93; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_94; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_95; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_96; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_97; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_98; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_99; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_100; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_101; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_102; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_103; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_104; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_105; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_106; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_107; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_108; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_109; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_110; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_111; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_112; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_113; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_114; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_115; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_116; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_117; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_118; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_119; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_120; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_121; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_122; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_123; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_124; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_125; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_126; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_127; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_128; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_129; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_130; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_131; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_132; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_133; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_134; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_135; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_136; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_137; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_138; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_139; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_140; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_141; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_142; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_143; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_144; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_145; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_146; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_147; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_148; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_149; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_150; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_151; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_152; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_153; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_154; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_155; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_156; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_157; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_158; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_159; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_160; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_161; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_162; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_163; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_164; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_165; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_166; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_167; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_168; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_169; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_170; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_171; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_172; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_173; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_174; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_175; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_176; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_177; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_178; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_179; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_180; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_181; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_182; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_183; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_184; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_185; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_186; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_187; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_188; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_189; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_190; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_191; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_192; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_193; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_194; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_195; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_196; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_197; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_198; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_199; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_200; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_201; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_202; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_203; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_204; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_205; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_206; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_207; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_208; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_209; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_210; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_211; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_212; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_213; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_214; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_215; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_216; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_217; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_218; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_219; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_220; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_221; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_222; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_223; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_224; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_225; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_226; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_227; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_228; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_229; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_230; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_231; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_232; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_233; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_234; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_235; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_236; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_237; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_238; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_239; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_240; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_241; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_242; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_243; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_244; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_245; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_246; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_247; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_248; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_249; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_250; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_251; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_252; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_253; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_254; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_255; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_256; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_257; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_258; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_259; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_260; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_261; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_262; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_263; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_264; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_265; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_266; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_267; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_268; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_269; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_270; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_271; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_272; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_273; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_274; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_275; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_276; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_277; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_278; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_279; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_280; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_281; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_282; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_283; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_284; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_285; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_286; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_287; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_288; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_289; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_290; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_291; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_292; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_293; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_294; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_295; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_296; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_297; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_298; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_299; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_300; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_301; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_302; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_303; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_304; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_305; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_306; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_307; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_308; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_309; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_310; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_311; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_312; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_313; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_314; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_315; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_316; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_317; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_318; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_319; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_320; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_321; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_322; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_323; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_324; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_325; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_326; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_327; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_328; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_329; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_330; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_331; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_332; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_333; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_334; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_335; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_336; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_337; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_338; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_339; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_340; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_341; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_342; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_343; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_344; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_345; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_346; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_347; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_348; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_349; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_350; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_351; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_352; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_353; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_354; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_355; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_356; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_357; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_358; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_359; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_360; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_361; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_362; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_363; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_364; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_365; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_366; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_367; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_368; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_369; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_370; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_371; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_372; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_373; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_374; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_375; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_376; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_377; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_378; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_379; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_380; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_381; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_382; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_383; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_384; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_385; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_386; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_387; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_388; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_389; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_390; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_391; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_392; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_393; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_394; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_395; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_396; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_397; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_398; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_399; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_400; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_401; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_402; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_403; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_404; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_405; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_406; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_407; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_408; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_409; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_410; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_411; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_412; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_413; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_414; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_415; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_416; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_417; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_418; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_419; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_420; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_421; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_422; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_423; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_424; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_425; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_426; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_427; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_428; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_429; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_430; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_431; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_432; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_433; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_434; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_435; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_436; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_437; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_438; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_439; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_440; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_441; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_442; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_443; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_444; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_445; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_446; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_447; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_448; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_449; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_450; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_451; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_452; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_453; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_454; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_455; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_456; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_457; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_458; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_459; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_460; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_461; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_462; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_463; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_464; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_465; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_466; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_467; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_468; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_469; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_470; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_471; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_472; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_473; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_474; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_475; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_476; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_477; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_478; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_479; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_480; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_481; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_482; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_483; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_484; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_485; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_486; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_487; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_488; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_489; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_490; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_491; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_492; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_493; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_494; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_495; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_496; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_497; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_498; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_499; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_500; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_501; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_502; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_503; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_504; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_505; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_506; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_507; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_508; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_509; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_510; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_511; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_512; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_513; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_514; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_515; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_516; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_517; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_518; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_519; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_520; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_521; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_522; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_523; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_524; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_525; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_526; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_527; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_528; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_529; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_530; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_531; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_532; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_533; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_534; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_535; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_536; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_537; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_538; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_539; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_540; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_541; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_542; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_543; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_544; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_545; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_546; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_547; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_548; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_549; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_550; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_551; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_552; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_553; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_554; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_555; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_556; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_557; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_558; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_559; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_560; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_561; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_562; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_563; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_564; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_565; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_566; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_567; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_568; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_569; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_570; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_571; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_572; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_573; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_574; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_575; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_576; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_577; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_578; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_579; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_580; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_581; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_582; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_583; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_584; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_585; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_586; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_587; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_588; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_589; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_590; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_591; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_592; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_593; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_594; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_595; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_596; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_597; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_598; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_599; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_600; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_601; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_602; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_603; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_604; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_605; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_606; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_607; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_608; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_609; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_610; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_611; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_612; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_613; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_614; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_615; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_616; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_617; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_618; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_619; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_620; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_621; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_622; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_623; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_624; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_625; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_626; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_627; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_628; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_629; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_630; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_631; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_632; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_633; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_634; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_635; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_636; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_637; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_638; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_639; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_640; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_641; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_642; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_643; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_644; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_645; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_646; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_647; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_648; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_649; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_650; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_651; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_652; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_653; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_654; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_655; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_656; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_657; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_658; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_659; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_660; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_661; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_662; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_663; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_664; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_665; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_666; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_667; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_668; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_669; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_670; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_671; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_672; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_673; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_674; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_675; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_676; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_677; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_678; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_679; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_680; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_681; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_682; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_683; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_684; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_685; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_686; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_687; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_688; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_689; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_690; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_691; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_692; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_693; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_694; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_695; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_696; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_697; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_698; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_699; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_700; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_701; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_702; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_703; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_704; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_705; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_706; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_707; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_708; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_709; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_710; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_711; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_712; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_713; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_714; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_715; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_716; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_717; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_718; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_719; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_720; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_721; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_722; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_723; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_724; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_725; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_726; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_727; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_728; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_729; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_730; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_731; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_732; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_733; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_734; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_735; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_736; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_737; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_738; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_739; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_740; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_741; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_742; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_743; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_744; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_745; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_746; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_747; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_748; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_749; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_750; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_751; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_752; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_753; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_754; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_755; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_756; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_757; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_758; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_759; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_760; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_761; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_762; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_763; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_764; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_765; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_766; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_767; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_768; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_769; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_770; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_771; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_772; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_773; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_774; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_775; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_776; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_777; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_778; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_779; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_780; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_781; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_782; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_783; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_784; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_785; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_786; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_787; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_788; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_789; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_790; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_791; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_792; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_793; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_794; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_795; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_796; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_797; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_798; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_799; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_800; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_801; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_802; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_803; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_804; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_805; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_806; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_807; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_808; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_809; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_810; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_811; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_812; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_813; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_814; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_815; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_816; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_817; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_818; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_819; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_820; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_821; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_822; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_823; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_824; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_825; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_826; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_827; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_828; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_829; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_830; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_831; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_832; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_833; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_834; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_835; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_836; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_837; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_838; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_839; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_840; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_841; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_842; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_843; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_844; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_845; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_846; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_847; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_848; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_849; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_850; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_851; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_852; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_853; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_854; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_855; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_856; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_857; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_858; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_859; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_860; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_861; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_862; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_863; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_864; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_865; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_866; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_867; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_868; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_869; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_870; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_871; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_872; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_873; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_874; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_875; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_876; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_877; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_878; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_879; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_880; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_881; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_882; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_883; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_884; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_885; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_886; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_887; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_888; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_889; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_890; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_891; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_892; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_893; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_894; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_895; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_896; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_897; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_898; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_899; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_900; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_901; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_902; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_903; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_904; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_905; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_906; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_907; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_908; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_909; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_910; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_911; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_912; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_913; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_914; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_915; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_916; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_917; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_918; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_919; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_920; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_921; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_922; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_923; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_924; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_925; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_926; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_927; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_928; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_929; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_930; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_931; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_932; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_933; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_934; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_935; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_936; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_937; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_938; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_939; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_940; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_941; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_942; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_943; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_944; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_945; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_946; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_947; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_948; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_949; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_950; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_951; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_952; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_953; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_954; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_955; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_956; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_957; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_958; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_959; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_960; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_961; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_962; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_963; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_964; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_965; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_966; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_967; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_968; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_969; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_970; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_971; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_972; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_973; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_974; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_975; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_976; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_977; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_978; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_979; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_980; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_981; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_982; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_983; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_984; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_985; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_986; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_987; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_988; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_989; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_990; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_991; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_992; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_993; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_994; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_995; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_996; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_997; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_998; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_999; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1000; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1001; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1002; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1003; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1004; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1005; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1006; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1007; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1008; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1009; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1010; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1011; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1012; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1013; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1014; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1015; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1016; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1017; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1018; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1019; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1020; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1021; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1022; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1023; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1024; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1025; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1026; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1027; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1028; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1029; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1030; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1031; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1032; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1033; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1034; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1035; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1036; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1037; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1038; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1039; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1040; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1041; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1042; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1043; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1044; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1045; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1046; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1047; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1048; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1049; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1050; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1051; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1052; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1053; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1054; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1055; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1056; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1057; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1058; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1059; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1060; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1061; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1062; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1063; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1064; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1065; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1066; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1067; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1068; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1069; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1070; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1071; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1072; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1073; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1074; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1075; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1076; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1077; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1078; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1079; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1080; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1081; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1082; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1083; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1084; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1085; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1086; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1087; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1088; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1089; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1090; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1091; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1092; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1093; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1094; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1095; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1096; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1097; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1098; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1099; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1100; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1101; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1102; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1103; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1104; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1105; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1106; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1107; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1108; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1109; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1110; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1111; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1112; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1113; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1114; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1115; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1116; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1117; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1118; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1119; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1120; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1121; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1122; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1123; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1124; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1125; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1126; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1127; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1128; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1129; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1130; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1131; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1132; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1133; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1134; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1135; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1136; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1137; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1138; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1139; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1140; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1141; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1142; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1143; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1144; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1145; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1146; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1147; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1148; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1149; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1150; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1151; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1152; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1153; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1154; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1155; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1156; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1157; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1158; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1159; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1160; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1161; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1162; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1163; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1164; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1165; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1166; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1167; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1168; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1169; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1170; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1171; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1172; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1173; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1174; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1175; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1176; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1177; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1178; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1179; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1180; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1181; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1182; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1183; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1184; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1185; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1186; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1187; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1188; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1189; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1190; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1191; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1192; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1193; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1194; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1195; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1196; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1197; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1198; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1199; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1200; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1201; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1202; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1203; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1204; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1205; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1206; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1207; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1208; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1209; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1210; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1211; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1212; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1213; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1214; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1215; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1216; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1217; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1218; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1219; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1220; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1221; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1222; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1223; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1224; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1225; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1226; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1227; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1228; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1229; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1230; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1231; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1232; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1233; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1234; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1235; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1236; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1237; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1238; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1239; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1240; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1241; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1242; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1243; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1244; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1245; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1246; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1247; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1248; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1249; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1250; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1251; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1252; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1253; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1254; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1255; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1256; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1257; // @[FloatingPointDesigns.scala 2274:23]
  reg [31:0] regs_1258; // @[FloatingPointDesigns.scala 2274:23]
  FP_reciprocal_newfpu FP_reciprocal_newfpu ( // @[FloatingPointDesigns.scala 2279:28]
    .clock(FP_reciprocal_newfpu_clock),
    .reset(FP_reciprocal_newfpu_reset),
    .io_in_en(FP_reciprocal_newfpu_io_in_en),
    .io_in_a(FP_reciprocal_newfpu_io_in_a),
    .io_out_s(FP_reciprocal_newfpu_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 2282:28]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_en(FP_multiplier_10ccs_io_in_en),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  assign io_out_s = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2286:14]
  assign FP_reciprocal_newfpu_clock = clock;
  assign FP_reciprocal_newfpu_reset = reset;
  assign FP_reciprocal_newfpu_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2280:22]
  assign FP_reciprocal_newfpu_io_in_a = io_in_b; // @[FloatingPointDesigns.scala 2281:21]
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2283:22]
  assign FP_multiplier_10ccs_io_in_a = regs_1258; // @[FloatingPointDesigns.scala 2284:21]
  assign FP_multiplier_10ccs_io_in_b = FP_reciprocal_newfpu_io_out_s; // @[FloatingPointDesigns.scala 2285:21]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_0 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_0 <= io_in_a; // @[FloatingPointDesigns.scala 2275:13]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1 <= regs_0; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_2 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_2 <= regs_1; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_3 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_3 <= regs_2; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_4 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_4 <= regs_3; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_5 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_5 <= regs_4; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_6 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_6 <= regs_5; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_7 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_7 <= regs_6; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_8 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_8 <= regs_7; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_9 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_9 <= regs_8; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_10 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_10 <= regs_9; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_11 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_11 <= regs_10; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_12 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_12 <= regs_11; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_13 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_13 <= regs_12; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_14 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_14 <= regs_13; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_15 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_15 <= regs_14; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_16 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_16 <= regs_15; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_17 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_17 <= regs_16; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_18 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_18 <= regs_17; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_19 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_19 <= regs_18; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_20 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_20 <= regs_19; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_21 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_21 <= regs_20; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_22 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_22 <= regs_21; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_23 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_23 <= regs_22; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_24 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_24 <= regs_23; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_25 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_25 <= regs_24; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_26 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_26 <= regs_25; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_27 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_27 <= regs_26; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_28 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_28 <= regs_27; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_29 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_29 <= regs_28; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_30 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_30 <= regs_29; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_31 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_31 <= regs_30; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_32 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_32 <= regs_31; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_33 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_33 <= regs_32; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_34 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_34 <= regs_33; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_35 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_35 <= regs_34; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_36 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_36 <= regs_35; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_37 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_37 <= regs_36; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_38 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_38 <= regs_37; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_39 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_39 <= regs_38; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_40 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_40 <= regs_39; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_41 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_41 <= regs_40; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_42 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_42 <= regs_41; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_43 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_43 <= regs_42; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_44 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_44 <= regs_43; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_45 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_45 <= regs_44; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_46 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_46 <= regs_45; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_47 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_47 <= regs_46; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_48 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_48 <= regs_47; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_49 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_49 <= regs_48; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_50 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_50 <= regs_49; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_51 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_51 <= regs_50; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_52 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_52 <= regs_51; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_53 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_53 <= regs_52; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_54 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_54 <= regs_53; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_55 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_55 <= regs_54; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_56 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_56 <= regs_55; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_57 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_57 <= regs_56; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_58 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_58 <= regs_57; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_59 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_59 <= regs_58; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_60 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_60 <= regs_59; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_61 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_61 <= regs_60; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_62 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_62 <= regs_61; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_63 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_63 <= regs_62; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_64 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_64 <= regs_63; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_65 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_65 <= regs_64; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_66 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_66 <= regs_65; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_67 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_67 <= regs_66; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_68 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_68 <= regs_67; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_69 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_69 <= regs_68; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_70 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_70 <= regs_69; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_71 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_71 <= regs_70; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_72 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_72 <= regs_71; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_73 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_73 <= regs_72; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_74 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_74 <= regs_73; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_75 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_75 <= regs_74; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_76 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_76 <= regs_75; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_77 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_77 <= regs_76; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_78 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_78 <= regs_77; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_79 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_79 <= regs_78; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_80 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_80 <= regs_79; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_81 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_81 <= regs_80; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_82 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_82 <= regs_81; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_83 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_83 <= regs_82; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_84 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_84 <= regs_83; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_85 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_85 <= regs_84; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_86 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_86 <= regs_85; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_87 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_87 <= regs_86; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_88 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_88 <= regs_87; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_89 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_89 <= regs_88; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_90 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_90 <= regs_89; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_91 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_91 <= regs_90; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_92 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_92 <= regs_91; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_93 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_93 <= regs_92; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_94 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_94 <= regs_93; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_95 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_95 <= regs_94; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_96 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_96 <= regs_95; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_97 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_97 <= regs_96; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_98 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_98 <= regs_97; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_99 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_99 <= regs_98; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_100 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_100 <= regs_99; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_101 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_101 <= regs_100; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_102 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_102 <= regs_101; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_103 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_103 <= regs_102; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_104 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_104 <= regs_103; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_105 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_105 <= regs_104; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_106 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_106 <= regs_105; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_107 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_107 <= regs_106; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_108 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_108 <= regs_107; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_109 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_109 <= regs_108; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_110 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_110 <= regs_109; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_111 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_111 <= regs_110; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_112 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_112 <= regs_111; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_113 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_113 <= regs_112; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_114 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_114 <= regs_113; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_115 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_115 <= regs_114; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_116 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_116 <= regs_115; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_117 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_117 <= regs_116; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_118 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_118 <= regs_117; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_119 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_119 <= regs_118; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_120 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_120 <= regs_119; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_121 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_121 <= regs_120; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_122 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_122 <= regs_121; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_123 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_123 <= regs_122; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_124 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_124 <= regs_123; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_125 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_125 <= regs_124; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_126 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_126 <= regs_125; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_127 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_127 <= regs_126; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_128 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_128 <= regs_127; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_129 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_129 <= regs_128; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_130 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_130 <= regs_129; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_131 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_131 <= regs_130; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_132 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_132 <= regs_131; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_133 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_133 <= regs_132; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_134 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_134 <= regs_133; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_135 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_135 <= regs_134; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_136 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_136 <= regs_135; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_137 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_137 <= regs_136; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_138 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_138 <= regs_137; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_139 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_139 <= regs_138; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_140 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_140 <= regs_139; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_141 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_141 <= regs_140; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_142 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_142 <= regs_141; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_143 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_143 <= regs_142; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_144 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_144 <= regs_143; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_145 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_145 <= regs_144; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_146 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_146 <= regs_145; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_147 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_147 <= regs_146; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_148 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_148 <= regs_147; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_149 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_149 <= regs_148; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_150 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_150 <= regs_149; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_151 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_151 <= regs_150; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_152 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_152 <= regs_151; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_153 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_153 <= regs_152; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_154 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_154 <= regs_153; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_155 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_155 <= regs_154; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_156 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_156 <= regs_155; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_157 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_157 <= regs_156; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_158 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_158 <= regs_157; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_159 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_159 <= regs_158; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_160 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_160 <= regs_159; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_161 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_161 <= regs_160; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_162 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_162 <= regs_161; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_163 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_163 <= regs_162; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_164 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_164 <= regs_163; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_165 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_165 <= regs_164; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_166 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_166 <= regs_165; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_167 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_167 <= regs_166; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_168 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_168 <= regs_167; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_169 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_169 <= regs_168; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_170 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_170 <= regs_169; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_171 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_171 <= regs_170; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_172 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_172 <= regs_171; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_173 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_173 <= regs_172; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_174 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_174 <= regs_173; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_175 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_175 <= regs_174; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_176 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_176 <= regs_175; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_177 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_177 <= regs_176; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_178 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_178 <= regs_177; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_179 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_179 <= regs_178; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_180 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_180 <= regs_179; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_181 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_181 <= regs_180; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_182 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_182 <= regs_181; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_183 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_183 <= regs_182; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_184 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_184 <= regs_183; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_185 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_185 <= regs_184; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_186 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_186 <= regs_185; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_187 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_187 <= regs_186; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_188 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_188 <= regs_187; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_189 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_189 <= regs_188; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_190 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_190 <= regs_189; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_191 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_191 <= regs_190; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_192 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_192 <= regs_191; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_193 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_193 <= regs_192; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_194 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_194 <= regs_193; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_195 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_195 <= regs_194; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_196 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_196 <= regs_195; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_197 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_197 <= regs_196; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_198 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_198 <= regs_197; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_199 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_199 <= regs_198; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_200 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_200 <= regs_199; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_201 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_201 <= regs_200; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_202 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_202 <= regs_201; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_203 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_203 <= regs_202; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_204 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_204 <= regs_203; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_205 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_205 <= regs_204; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_206 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_206 <= regs_205; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_207 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_207 <= regs_206; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_208 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_208 <= regs_207; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_209 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_209 <= regs_208; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_210 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_210 <= regs_209; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_211 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_211 <= regs_210; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_212 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_212 <= regs_211; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_213 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_213 <= regs_212; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_214 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_214 <= regs_213; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_215 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_215 <= regs_214; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_216 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_216 <= regs_215; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_217 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_217 <= regs_216; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_218 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_218 <= regs_217; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_219 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_219 <= regs_218; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_220 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_220 <= regs_219; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_221 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_221 <= regs_220; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_222 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_222 <= regs_221; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_223 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_223 <= regs_222; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_224 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_224 <= regs_223; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_225 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_225 <= regs_224; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_226 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_226 <= regs_225; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_227 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_227 <= regs_226; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_228 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_228 <= regs_227; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_229 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_229 <= regs_228; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_230 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_230 <= regs_229; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_231 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_231 <= regs_230; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_232 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_232 <= regs_231; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_233 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_233 <= regs_232; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_234 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_234 <= regs_233; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_235 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_235 <= regs_234; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_236 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_236 <= regs_235; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_237 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_237 <= regs_236; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_238 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_238 <= regs_237; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_239 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_239 <= regs_238; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_240 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_240 <= regs_239; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_241 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_241 <= regs_240; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_242 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_242 <= regs_241; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_243 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_243 <= regs_242; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_244 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_244 <= regs_243; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_245 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_245 <= regs_244; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_246 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_246 <= regs_245; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_247 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_247 <= regs_246; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_248 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_248 <= regs_247; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_249 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_249 <= regs_248; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_250 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_250 <= regs_249; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_251 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_251 <= regs_250; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_252 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_252 <= regs_251; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_253 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_253 <= regs_252; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_254 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_254 <= regs_253; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_255 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_255 <= regs_254; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_256 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_256 <= regs_255; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_257 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_257 <= regs_256; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_258 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_258 <= regs_257; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_259 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_259 <= regs_258; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_260 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_260 <= regs_259; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_261 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_261 <= regs_260; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_262 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_262 <= regs_261; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_263 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_263 <= regs_262; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_264 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_264 <= regs_263; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_265 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_265 <= regs_264; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_266 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_266 <= regs_265; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_267 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_267 <= regs_266; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_268 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_268 <= regs_267; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_269 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_269 <= regs_268; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_270 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_270 <= regs_269; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_271 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_271 <= regs_270; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_272 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_272 <= regs_271; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_273 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_273 <= regs_272; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_274 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_274 <= regs_273; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_275 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_275 <= regs_274; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_276 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_276 <= regs_275; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_277 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_277 <= regs_276; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_278 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_278 <= regs_277; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_279 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_279 <= regs_278; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_280 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_280 <= regs_279; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_281 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_281 <= regs_280; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_282 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_282 <= regs_281; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_283 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_283 <= regs_282; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_284 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_284 <= regs_283; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_285 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_285 <= regs_284; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_286 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_286 <= regs_285; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_287 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_287 <= regs_286; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_288 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_288 <= regs_287; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_289 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_289 <= regs_288; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_290 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_290 <= regs_289; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_291 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_291 <= regs_290; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_292 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_292 <= regs_291; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_293 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_293 <= regs_292; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_294 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_294 <= regs_293; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_295 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_295 <= regs_294; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_296 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_296 <= regs_295; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_297 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_297 <= regs_296; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_298 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_298 <= regs_297; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_299 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_299 <= regs_298; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_300 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_300 <= regs_299; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_301 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_301 <= regs_300; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_302 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_302 <= regs_301; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_303 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_303 <= regs_302; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_304 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_304 <= regs_303; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_305 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_305 <= regs_304; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_306 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_306 <= regs_305; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_307 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_307 <= regs_306; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_308 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_308 <= regs_307; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_309 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_309 <= regs_308; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_310 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_310 <= regs_309; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_311 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_311 <= regs_310; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_312 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_312 <= regs_311; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_313 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_313 <= regs_312; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_314 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_314 <= regs_313; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_315 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_315 <= regs_314; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_316 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_316 <= regs_315; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_317 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_317 <= regs_316; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_318 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_318 <= regs_317; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_319 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_319 <= regs_318; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_320 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_320 <= regs_319; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_321 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_321 <= regs_320; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_322 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_322 <= regs_321; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_323 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_323 <= regs_322; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_324 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_324 <= regs_323; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_325 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_325 <= regs_324; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_326 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_326 <= regs_325; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_327 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_327 <= regs_326; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_328 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_328 <= regs_327; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_329 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_329 <= regs_328; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_330 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_330 <= regs_329; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_331 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_331 <= regs_330; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_332 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_332 <= regs_331; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_333 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_333 <= regs_332; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_334 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_334 <= regs_333; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_335 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_335 <= regs_334; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_336 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_336 <= regs_335; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_337 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_337 <= regs_336; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_338 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_338 <= regs_337; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_339 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_339 <= regs_338; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_340 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_340 <= regs_339; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_341 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_341 <= regs_340; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_342 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_342 <= regs_341; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_343 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_343 <= regs_342; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_344 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_344 <= regs_343; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_345 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_345 <= regs_344; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_346 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_346 <= regs_345; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_347 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_347 <= regs_346; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_348 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_348 <= regs_347; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_349 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_349 <= regs_348; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_350 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_350 <= regs_349; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_351 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_351 <= regs_350; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_352 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_352 <= regs_351; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_353 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_353 <= regs_352; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_354 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_354 <= regs_353; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_355 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_355 <= regs_354; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_356 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_356 <= regs_355; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_357 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_357 <= regs_356; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_358 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_358 <= regs_357; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_359 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_359 <= regs_358; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_360 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_360 <= regs_359; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_361 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_361 <= regs_360; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_362 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_362 <= regs_361; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_363 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_363 <= regs_362; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_364 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_364 <= regs_363; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_365 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_365 <= regs_364; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_366 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_366 <= regs_365; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_367 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_367 <= regs_366; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_368 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_368 <= regs_367; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_369 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_369 <= regs_368; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_370 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_370 <= regs_369; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_371 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_371 <= regs_370; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_372 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_372 <= regs_371; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_373 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_373 <= regs_372; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_374 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_374 <= regs_373; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_375 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_375 <= regs_374; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_376 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_376 <= regs_375; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_377 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_377 <= regs_376; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_378 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_378 <= regs_377; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_379 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_379 <= regs_378; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_380 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_380 <= regs_379; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_381 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_381 <= regs_380; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_382 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_382 <= regs_381; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_383 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_383 <= regs_382; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_384 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_384 <= regs_383; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_385 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_385 <= regs_384; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_386 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_386 <= regs_385; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_387 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_387 <= regs_386; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_388 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_388 <= regs_387; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_389 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_389 <= regs_388; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_390 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_390 <= regs_389; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_391 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_391 <= regs_390; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_392 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_392 <= regs_391; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_393 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_393 <= regs_392; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_394 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_394 <= regs_393; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_395 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_395 <= regs_394; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_396 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_396 <= regs_395; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_397 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_397 <= regs_396; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_398 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_398 <= regs_397; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_399 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_399 <= regs_398; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_400 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_400 <= regs_399; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_401 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_401 <= regs_400; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_402 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_402 <= regs_401; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_403 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_403 <= regs_402; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_404 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_404 <= regs_403; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_405 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_405 <= regs_404; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_406 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_406 <= regs_405; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_407 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_407 <= regs_406; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_408 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_408 <= regs_407; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_409 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_409 <= regs_408; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_410 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_410 <= regs_409; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_411 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_411 <= regs_410; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_412 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_412 <= regs_411; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_413 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_413 <= regs_412; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_414 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_414 <= regs_413; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_415 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_415 <= regs_414; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_416 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_416 <= regs_415; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_417 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_417 <= regs_416; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_418 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_418 <= regs_417; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_419 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_419 <= regs_418; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_420 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_420 <= regs_419; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_421 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_421 <= regs_420; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_422 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_422 <= regs_421; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_423 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_423 <= regs_422; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_424 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_424 <= regs_423; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_425 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_425 <= regs_424; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_426 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_426 <= regs_425; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_427 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_427 <= regs_426; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_428 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_428 <= regs_427; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_429 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_429 <= regs_428; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_430 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_430 <= regs_429; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_431 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_431 <= regs_430; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_432 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_432 <= regs_431; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_433 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_433 <= regs_432; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_434 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_434 <= regs_433; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_435 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_435 <= regs_434; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_436 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_436 <= regs_435; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_437 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_437 <= regs_436; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_438 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_438 <= regs_437; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_439 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_439 <= regs_438; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_440 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_440 <= regs_439; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_441 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_441 <= regs_440; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_442 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_442 <= regs_441; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_443 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_443 <= regs_442; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_444 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_444 <= regs_443; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_445 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_445 <= regs_444; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_446 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_446 <= regs_445; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_447 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_447 <= regs_446; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_448 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_448 <= regs_447; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_449 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_449 <= regs_448; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_450 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_450 <= regs_449; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_451 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_451 <= regs_450; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_452 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_452 <= regs_451; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_453 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_453 <= regs_452; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_454 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_454 <= regs_453; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_455 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_455 <= regs_454; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_456 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_456 <= regs_455; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_457 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_457 <= regs_456; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_458 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_458 <= regs_457; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_459 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_459 <= regs_458; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_460 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_460 <= regs_459; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_461 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_461 <= regs_460; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_462 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_462 <= regs_461; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_463 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_463 <= regs_462; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_464 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_464 <= regs_463; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_465 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_465 <= regs_464; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_466 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_466 <= regs_465; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_467 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_467 <= regs_466; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_468 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_468 <= regs_467; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_469 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_469 <= regs_468; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_470 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_470 <= regs_469; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_471 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_471 <= regs_470; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_472 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_472 <= regs_471; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_473 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_473 <= regs_472; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_474 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_474 <= regs_473; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_475 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_475 <= regs_474; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_476 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_476 <= regs_475; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_477 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_477 <= regs_476; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_478 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_478 <= regs_477; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_479 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_479 <= regs_478; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_480 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_480 <= regs_479; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_481 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_481 <= regs_480; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_482 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_482 <= regs_481; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_483 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_483 <= regs_482; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_484 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_484 <= regs_483; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_485 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_485 <= regs_484; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_486 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_486 <= regs_485; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_487 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_487 <= regs_486; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_488 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_488 <= regs_487; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_489 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_489 <= regs_488; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_490 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_490 <= regs_489; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_491 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_491 <= regs_490; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_492 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_492 <= regs_491; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_493 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_493 <= regs_492; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_494 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_494 <= regs_493; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_495 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_495 <= regs_494; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_496 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_496 <= regs_495; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_497 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_497 <= regs_496; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_498 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_498 <= regs_497; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_499 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_499 <= regs_498; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_500 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_500 <= regs_499; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_501 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_501 <= regs_500; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_502 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_502 <= regs_501; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_503 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_503 <= regs_502; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_504 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_504 <= regs_503; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_505 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_505 <= regs_504; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_506 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_506 <= regs_505; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_507 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_507 <= regs_506; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_508 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_508 <= regs_507; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_509 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_509 <= regs_508; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_510 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_510 <= regs_509; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_511 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_511 <= regs_510; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_512 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_512 <= regs_511; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_513 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_513 <= regs_512; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_514 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_514 <= regs_513; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_515 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_515 <= regs_514; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_516 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_516 <= regs_515; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_517 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_517 <= regs_516; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_518 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_518 <= regs_517; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_519 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_519 <= regs_518; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_520 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_520 <= regs_519; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_521 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_521 <= regs_520; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_522 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_522 <= regs_521; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_523 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_523 <= regs_522; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_524 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_524 <= regs_523; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_525 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_525 <= regs_524; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_526 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_526 <= regs_525; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_527 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_527 <= regs_526; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_528 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_528 <= regs_527; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_529 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_529 <= regs_528; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_530 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_530 <= regs_529; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_531 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_531 <= regs_530; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_532 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_532 <= regs_531; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_533 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_533 <= regs_532; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_534 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_534 <= regs_533; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_535 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_535 <= regs_534; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_536 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_536 <= regs_535; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_537 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_537 <= regs_536; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_538 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_538 <= regs_537; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_539 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_539 <= regs_538; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_540 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_540 <= regs_539; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_541 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_541 <= regs_540; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_542 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_542 <= regs_541; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_543 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_543 <= regs_542; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_544 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_544 <= regs_543; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_545 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_545 <= regs_544; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_546 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_546 <= regs_545; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_547 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_547 <= regs_546; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_548 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_548 <= regs_547; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_549 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_549 <= regs_548; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_550 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_550 <= regs_549; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_551 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_551 <= regs_550; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_552 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_552 <= regs_551; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_553 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_553 <= regs_552; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_554 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_554 <= regs_553; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_555 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_555 <= regs_554; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_556 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_556 <= regs_555; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_557 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_557 <= regs_556; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_558 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_558 <= regs_557; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_559 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_559 <= regs_558; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_560 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_560 <= regs_559; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_561 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_561 <= regs_560; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_562 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_562 <= regs_561; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_563 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_563 <= regs_562; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_564 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_564 <= regs_563; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_565 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_565 <= regs_564; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_566 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_566 <= regs_565; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_567 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_567 <= regs_566; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_568 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_568 <= regs_567; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_569 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_569 <= regs_568; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_570 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_570 <= regs_569; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_571 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_571 <= regs_570; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_572 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_572 <= regs_571; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_573 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_573 <= regs_572; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_574 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_574 <= regs_573; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_575 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_575 <= regs_574; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_576 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_576 <= regs_575; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_577 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_577 <= regs_576; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_578 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_578 <= regs_577; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_579 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_579 <= regs_578; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_580 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_580 <= regs_579; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_581 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_581 <= regs_580; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_582 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_582 <= regs_581; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_583 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_583 <= regs_582; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_584 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_584 <= regs_583; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_585 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_585 <= regs_584; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_586 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_586 <= regs_585; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_587 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_587 <= regs_586; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_588 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_588 <= regs_587; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_589 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_589 <= regs_588; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_590 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_590 <= regs_589; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_591 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_591 <= regs_590; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_592 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_592 <= regs_591; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_593 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_593 <= regs_592; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_594 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_594 <= regs_593; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_595 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_595 <= regs_594; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_596 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_596 <= regs_595; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_597 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_597 <= regs_596; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_598 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_598 <= regs_597; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_599 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_599 <= regs_598; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_600 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_600 <= regs_599; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_601 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_601 <= regs_600; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_602 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_602 <= regs_601; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_603 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_603 <= regs_602; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_604 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_604 <= regs_603; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_605 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_605 <= regs_604; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_606 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_606 <= regs_605; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_607 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_607 <= regs_606; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_608 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_608 <= regs_607; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_609 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_609 <= regs_608; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_610 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_610 <= regs_609; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_611 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_611 <= regs_610; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_612 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_612 <= regs_611; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_613 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_613 <= regs_612; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_614 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_614 <= regs_613; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_615 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_615 <= regs_614; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_616 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_616 <= regs_615; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_617 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_617 <= regs_616; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_618 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_618 <= regs_617; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_619 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_619 <= regs_618; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_620 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_620 <= regs_619; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_621 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_621 <= regs_620; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_622 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_622 <= regs_621; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_623 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_623 <= regs_622; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_624 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_624 <= regs_623; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_625 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_625 <= regs_624; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_626 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_626 <= regs_625; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_627 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_627 <= regs_626; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_628 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_628 <= regs_627; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_629 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_629 <= regs_628; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_630 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_630 <= regs_629; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_631 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_631 <= regs_630; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_632 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_632 <= regs_631; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_633 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_633 <= regs_632; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_634 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_634 <= regs_633; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_635 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_635 <= regs_634; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_636 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_636 <= regs_635; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_637 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_637 <= regs_636; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_638 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_638 <= regs_637; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_639 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_639 <= regs_638; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_640 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_640 <= regs_639; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_641 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_641 <= regs_640; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_642 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_642 <= regs_641; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_643 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_643 <= regs_642; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_644 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_644 <= regs_643; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_645 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_645 <= regs_644; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_646 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_646 <= regs_645; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_647 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_647 <= regs_646; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_648 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_648 <= regs_647; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_649 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_649 <= regs_648; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_650 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_650 <= regs_649; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_651 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_651 <= regs_650; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_652 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_652 <= regs_651; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_653 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_653 <= regs_652; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_654 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_654 <= regs_653; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_655 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_655 <= regs_654; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_656 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_656 <= regs_655; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_657 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_657 <= regs_656; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_658 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_658 <= regs_657; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_659 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_659 <= regs_658; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_660 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_660 <= regs_659; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_661 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_661 <= regs_660; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_662 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_662 <= regs_661; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_663 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_663 <= regs_662; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_664 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_664 <= regs_663; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_665 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_665 <= regs_664; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_666 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_666 <= regs_665; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_667 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_667 <= regs_666; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_668 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_668 <= regs_667; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_669 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_669 <= regs_668; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_670 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_670 <= regs_669; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_671 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_671 <= regs_670; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_672 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_672 <= regs_671; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_673 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_673 <= regs_672; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_674 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_674 <= regs_673; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_675 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_675 <= regs_674; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_676 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_676 <= regs_675; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_677 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_677 <= regs_676; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_678 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_678 <= regs_677; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_679 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_679 <= regs_678; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_680 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_680 <= regs_679; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_681 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_681 <= regs_680; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_682 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_682 <= regs_681; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_683 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_683 <= regs_682; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_684 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_684 <= regs_683; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_685 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_685 <= regs_684; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_686 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_686 <= regs_685; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_687 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_687 <= regs_686; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_688 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_688 <= regs_687; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_689 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_689 <= regs_688; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_690 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_690 <= regs_689; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_691 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_691 <= regs_690; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_692 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_692 <= regs_691; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_693 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_693 <= regs_692; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_694 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_694 <= regs_693; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_695 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_695 <= regs_694; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_696 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_696 <= regs_695; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_697 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_697 <= regs_696; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_698 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_698 <= regs_697; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_699 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_699 <= regs_698; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_700 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_700 <= regs_699; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_701 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_701 <= regs_700; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_702 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_702 <= regs_701; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_703 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_703 <= regs_702; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_704 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_704 <= regs_703; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_705 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_705 <= regs_704; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_706 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_706 <= regs_705; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_707 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_707 <= regs_706; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_708 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_708 <= regs_707; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_709 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_709 <= regs_708; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_710 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_710 <= regs_709; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_711 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_711 <= regs_710; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_712 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_712 <= regs_711; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_713 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_713 <= regs_712; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_714 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_714 <= regs_713; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_715 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_715 <= regs_714; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_716 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_716 <= regs_715; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_717 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_717 <= regs_716; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_718 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_718 <= regs_717; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_719 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_719 <= regs_718; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_720 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_720 <= regs_719; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_721 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_721 <= regs_720; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_722 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_722 <= regs_721; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_723 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_723 <= regs_722; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_724 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_724 <= regs_723; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_725 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_725 <= regs_724; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_726 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_726 <= regs_725; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_727 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_727 <= regs_726; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_728 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_728 <= regs_727; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_729 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_729 <= regs_728; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_730 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_730 <= regs_729; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_731 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_731 <= regs_730; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_732 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_732 <= regs_731; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_733 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_733 <= regs_732; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_734 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_734 <= regs_733; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_735 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_735 <= regs_734; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_736 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_736 <= regs_735; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_737 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_737 <= regs_736; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_738 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_738 <= regs_737; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_739 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_739 <= regs_738; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_740 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_740 <= regs_739; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_741 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_741 <= regs_740; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_742 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_742 <= regs_741; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_743 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_743 <= regs_742; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_744 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_744 <= regs_743; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_745 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_745 <= regs_744; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_746 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_746 <= regs_745; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_747 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_747 <= regs_746; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_748 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_748 <= regs_747; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_749 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_749 <= regs_748; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_750 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_750 <= regs_749; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_751 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_751 <= regs_750; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_752 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_752 <= regs_751; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_753 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_753 <= regs_752; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_754 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_754 <= regs_753; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_755 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_755 <= regs_754; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_756 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_756 <= regs_755; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_757 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_757 <= regs_756; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_758 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_758 <= regs_757; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_759 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_759 <= regs_758; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_760 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_760 <= regs_759; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_761 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_761 <= regs_760; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_762 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_762 <= regs_761; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_763 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_763 <= regs_762; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_764 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_764 <= regs_763; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_765 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_765 <= regs_764; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_766 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_766 <= regs_765; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_767 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_767 <= regs_766; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_768 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_768 <= regs_767; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_769 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_769 <= regs_768; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_770 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_770 <= regs_769; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_771 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_771 <= regs_770; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_772 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_772 <= regs_771; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_773 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_773 <= regs_772; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_774 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_774 <= regs_773; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_775 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_775 <= regs_774; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_776 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_776 <= regs_775; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_777 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_777 <= regs_776; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_778 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_778 <= regs_777; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_779 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_779 <= regs_778; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_780 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_780 <= regs_779; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_781 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_781 <= regs_780; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_782 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_782 <= regs_781; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_783 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_783 <= regs_782; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_784 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_784 <= regs_783; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_785 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_785 <= regs_784; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_786 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_786 <= regs_785; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_787 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_787 <= regs_786; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_788 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_788 <= regs_787; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_789 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_789 <= regs_788; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_790 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_790 <= regs_789; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_791 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_791 <= regs_790; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_792 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_792 <= regs_791; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_793 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_793 <= regs_792; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_794 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_794 <= regs_793; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_795 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_795 <= regs_794; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_796 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_796 <= regs_795; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_797 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_797 <= regs_796; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_798 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_798 <= regs_797; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_799 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_799 <= regs_798; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_800 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_800 <= regs_799; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_801 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_801 <= regs_800; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_802 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_802 <= regs_801; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_803 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_803 <= regs_802; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_804 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_804 <= regs_803; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_805 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_805 <= regs_804; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_806 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_806 <= regs_805; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_807 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_807 <= regs_806; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_808 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_808 <= regs_807; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_809 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_809 <= regs_808; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_810 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_810 <= regs_809; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_811 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_811 <= regs_810; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_812 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_812 <= regs_811; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_813 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_813 <= regs_812; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_814 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_814 <= regs_813; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_815 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_815 <= regs_814; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_816 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_816 <= regs_815; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_817 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_817 <= regs_816; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_818 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_818 <= regs_817; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_819 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_819 <= regs_818; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_820 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_820 <= regs_819; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_821 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_821 <= regs_820; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_822 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_822 <= regs_821; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_823 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_823 <= regs_822; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_824 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_824 <= regs_823; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_825 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_825 <= regs_824; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_826 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_826 <= regs_825; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_827 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_827 <= regs_826; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_828 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_828 <= regs_827; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_829 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_829 <= regs_828; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_830 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_830 <= regs_829; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_831 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_831 <= regs_830; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_832 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_832 <= regs_831; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_833 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_833 <= regs_832; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_834 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_834 <= regs_833; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_835 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_835 <= regs_834; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_836 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_836 <= regs_835; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_837 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_837 <= regs_836; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_838 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_838 <= regs_837; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_839 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_839 <= regs_838; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_840 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_840 <= regs_839; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_841 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_841 <= regs_840; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_842 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_842 <= regs_841; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_843 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_843 <= regs_842; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_844 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_844 <= regs_843; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_845 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_845 <= regs_844; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_846 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_846 <= regs_845; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_847 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_847 <= regs_846; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_848 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_848 <= regs_847; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_849 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_849 <= regs_848; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_850 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_850 <= regs_849; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_851 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_851 <= regs_850; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_852 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_852 <= regs_851; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_853 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_853 <= regs_852; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_854 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_854 <= regs_853; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_855 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_855 <= regs_854; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_856 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_856 <= regs_855; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_857 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_857 <= regs_856; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_858 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_858 <= regs_857; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_859 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_859 <= regs_858; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_860 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_860 <= regs_859; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_861 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_861 <= regs_860; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_862 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_862 <= regs_861; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_863 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_863 <= regs_862; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_864 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_864 <= regs_863; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_865 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_865 <= regs_864; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_866 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_866 <= regs_865; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_867 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_867 <= regs_866; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_868 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_868 <= regs_867; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_869 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_869 <= regs_868; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_870 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_870 <= regs_869; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_871 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_871 <= regs_870; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_872 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_872 <= regs_871; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_873 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_873 <= regs_872; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_874 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_874 <= regs_873; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_875 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_875 <= regs_874; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_876 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_876 <= regs_875; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_877 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_877 <= regs_876; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_878 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_878 <= regs_877; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_879 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_879 <= regs_878; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_880 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_880 <= regs_879; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_881 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_881 <= regs_880; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_882 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_882 <= regs_881; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_883 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_883 <= regs_882; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_884 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_884 <= regs_883; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_885 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_885 <= regs_884; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_886 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_886 <= regs_885; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_887 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_887 <= regs_886; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_888 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_888 <= regs_887; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_889 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_889 <= regs_888; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_890 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_890 <= regs_889; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_891 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_891 <= regs_890; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_892 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_892 <= regs_891; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_893 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_893 <= regs_892; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_894 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_894 <= regs_893; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_895 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_895 <= regs_894; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_896 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_896 <= regs_895; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_897 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_897 <= regs_896; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_898 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_898 <= regs_897; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_899 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_899 <= regs_898; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_900 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_900 <= regs_899; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_901 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_901 <= regs_900; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_902 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_902 <= regs_901; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_903 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_903 <= regs_902; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_904 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_904 <= regs_903; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_905 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_905 <= regs_904; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_906 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_906 <= regs_905; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_907 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_907 <= regs_906; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_908 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_908 <= regs_907; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_909 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_909 <= regs_908; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_910 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_910 <= regs_909; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_911 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_911 <= regs_910; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_912 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_912 <= regs_911; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_913 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_913 <= regs_912; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_914 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_914 <= regs_913; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_915 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_915 <= regs_914; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_916 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_916 <= regs_915; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_917 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_917 <= regs_916; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_918 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_918 <= regs_917; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_919 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_919 <= regs_918; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_920 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_920 <= regs_919; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_921 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_921 <= regs_920; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_922 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_922 <= regs_921; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_923 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_923 <= regs_922; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_924 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_924 <= regs_923; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_925 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_925 <= regs_924; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_926 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_926 <= regs_925; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_927 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_927 <= regs_926; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_928 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_928 <= regs_927; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_929 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_929 <= regs_928; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_930 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_930 <= regs_929; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_931 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_931 <= regs_930; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_932 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_932 <= regs_931; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_933 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_933 <= regs_932; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_934 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_934 <= regs_933; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_935 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_935 <= regs_934; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_936 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_936 <= regs_935; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_937 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_937 <= regs_936; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_938 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_938 <= regs_937; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_939 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_939 <= regs_938; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_940 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_940 <= regs_939; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_941 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_941 <= regs_940; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_942 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_942 <= regs_941; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_943 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_943 <= regs_942; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_944 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_944 <= regs_943; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_945 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_945 <= regs_944; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_946 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_946 <= regs_945; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_947 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_947 <= regs_946; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_948 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_948 <= regs_947; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_949 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_949 <= regs_948; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_950 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_950 <= regs_949; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_951 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_951 <= regs_950; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_952 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_952 <= regs_951; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_953 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_953 <= regs_952; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_954 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_954 <= regs_953; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_955 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_955 <= regs_954; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_956 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_956 <= regs_955; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_957 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_957 <= regs_956; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_958 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_958 <= regs_957; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_959 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_959 <= regs_958; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_960 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_960 <= regs_959; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_961 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_961 <= regs_960; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_962 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_962 <= regs_961; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_963 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_963 <= regs_962; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_964 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_964 <= regs_963; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_965 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_965 <= regs_964; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_966 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_966 <= regs_965; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_967 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_967 <= regs_966; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_968 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_968 <= regs_967; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_969 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_969 <= regs_968; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_970 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_970 <= regs_969; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_971 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_971 <= regs_970; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_972 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_972 <= regs_971; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_973 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_973 <= regs_972; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_974 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_974 <= regs_973; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_975 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_975 <= regs_974; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_976 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_976 <= regs_975; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_977 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_977 <= regs_976; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_978 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_978 <= regs_977; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_979 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_979 <= regs_978; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_980 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_980 <= regs_979; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_981 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_981 <= regs_980; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_982 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_982 <= regs_981; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_983 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_983 <= regs_982; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_984 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_984 <= regs_983; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_985 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_985 <= regs_984; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_986 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_986 <= regs_985; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_987 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_987 <= regs_986; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_988 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_988 <= regs_987; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_989 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_989 <= regs_988; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_990 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_990 <= regs_989; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_991 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_991 <= regs_990; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_992 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_992 <= regs_991; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_993 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_993 <= regs_992; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_994 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_994 <= regs_993; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_995 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_995 <= regs_994; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_996 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_996 <= regs_995; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_997 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_997 <= regs_996; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_998 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_998 <= regs_997; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_999 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_999 <= regs_998; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1000 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1000 <= regs_999; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1001 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1001 <= regs_1000; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1002 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1002 <= regs_1001; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1003 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1003 <= regs_1002; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1004 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1004 <= regs_1003; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1005 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1005 <= regs_1004; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1006 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1006 <= regs_1005; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1007 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1007 <= regs_1006; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1008 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1008 <= regs_1007; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1009 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1009 <= regs_1008; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1010 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1010 <= regs_1009; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1011 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1011 <= regs_1010; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1012 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1012 <= regs_1011; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1013 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1013 <= regs_1012; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1014 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1014 <= regs_1013; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1015 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1015 <= regs_1014; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1016 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1016 <= regs_1015; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1017 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1017 <= regs_1016; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1018 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1018 <= regs_1017; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1019 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1019 <= regs_1018; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1020 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1020 <= regs_1019; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1021 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1021 <= regs_1020; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1022 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1022 <= regs_1021; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1023 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1023 <= regs_1022; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1024 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1024 <= regs_1023; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1025 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1025 <= regs_1024; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1026 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1026 <= regs_1025; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1027 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1027 <= regs_1026; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1028 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1028 <= regs_1027; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1029 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1029 <= regs_1028; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1030 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1030 <= regs_1029; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1031 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1031 <= regs_1030; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1032 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1032 <= regs_1031; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1033 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1033 <= regs_1032; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1034 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1034 <= regs_1033; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1035 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1035 <= regs_1034; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1036 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1036 <= regs_1035; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1037 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1037 <= regs_1036; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1038 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1038 <= regs_1037; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1039 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1039 <= regs_1038; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1040 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1040 <= regs_1039; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1041 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1041 <= regs_1040; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1042 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1042 <= regs_1041; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1043 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1043 <= regs_1042; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1044 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1044 <= regs_1043; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1045 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1045 <= regs_1044; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1046 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1046 <= regs_1045; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1047 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1047 <= regs_1046; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1048 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1048 <= regs_1047; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1049 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1049 <= regs_1048; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1050 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1050 <= regs_1049; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1051 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1051 <= regs_1050; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1052 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1052 <= regs_1051; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1053 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1053 <= regs_1052; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1054 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1054 <= regs_1053; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1055 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1055 <= regs_1054; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1056 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1056 <= regs_1055; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1057 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1057 <= regs_1056; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1058 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1058 <= regs_1057; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1059 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1059 <= regs_1058; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1060 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1060 <= regs_1059; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1061 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1061 <= regs_1060; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1062 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1062 <= regs_1061; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1063 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1063 <= regs_1062; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1064 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1064 <= regs_1063; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1065 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1065 <= regs_1064; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1066 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1066 <= regs_1065; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1067 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1067 <= regs_1066; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1068 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1068 <= regs_1067; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1069 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1069 <= regs_1068; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1070 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1070 <= regs_1069; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1071 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1071 <= regs_1070; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1072 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1072 <= regs_1071; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1073 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1073 <= regs_1072; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1074 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1074 <= regs_1073; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1075 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1075 <= regs_1074; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1076 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1076 <= regs_1075; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1077 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1077 <= regs_1076; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1078 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1078 <= regs_1077; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1079 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1079 <= regs_1078; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1080 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1080 <= regs_1079; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1081 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1081 <= regs_1080; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1082 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1082 <= regs_1081; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1083 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1083 <= regs_1082; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1084 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1084 <= regs_1083; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1085 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1085 <= regs_1084; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1086 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1086 <= regs_1085; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1087 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1087 <= regs_1086; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1088 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1088 <= regs_1087; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1089 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1089 <= regs_1088; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1090 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1090 <= regs_1089; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1091 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1091 <= regs_1090; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1092 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1092 <= regs_1091; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1093 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1093 <= regs_1092; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1094 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1094 <= regs_1093; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1095 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1095 <= regs_1094; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1096 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1096 <= regs_1095; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1097 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1097 <= regs_1096; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1098 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1098 <= regs_1097; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1099 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1099 <= regs_1098; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1100 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1100 <= regs_1099; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1101 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1101 <= regs_1100; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1102 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1102 <= regs_1101; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1103 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1103 <= regs_1102; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1104 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1104 <= regs_1103; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1105 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1105 <= regs_1104; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1106 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1106 <= regs_1105; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1107 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1107 <= regs_1106; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1108 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1108 <= regs_1107; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1109 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1109 <= regs_1108; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1110 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1110 <= regs_1109; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1111 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1111 <= regs_1110; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1112 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1112 <= regs_1111; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1113 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1113 <= regs_1112; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1114 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1114 <= regs_1113; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1115 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1115 <= regs_1114; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1116 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1116 <= regs_1115; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1117 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1117 <= regs_1116; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1118 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1118 <= regs_1117; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1119 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1119 <= regs_1118; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1120 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1120 <= regs_1119; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1121 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1121 <= regs_1120; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1122 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1122 <= regs_1121; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1123 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1123 <= regs_1122; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1124 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1124 <= regs_1123; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1125 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1125 <= regs_1124; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1126 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1126 <= regs_1125; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1127 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1127 <= regs_1126; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1128 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1128 <= regs_1127; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1129 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1129 <= regs_1128; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1130 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1130 <= regs_1129; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1131 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1131 <= regs_1130; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1132 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1132 <= regs_1131; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1133 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1133 <= regs_1132; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1134 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1134 <= regs_1133; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1135 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1135 <= regs_1134; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1136 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1136 <= regs_1135; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1137 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1137 <= regs_1136; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1138 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1138 <= regs_1137; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1139 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1139 <= regs_1138; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1140 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1140 <= regs_1139; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1141 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1141 <= regs_1140; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1142 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1142 <= regs_1141; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1143 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1143 <= regs_1142; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1144 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1144 <= regs_1143; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1145 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1145 <= regs_1144; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1146 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1146 <= regs_1145; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1147 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1147 <= regs_1146; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1148 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1148 <= regs_1147; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1149 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1149 <= regs_1148; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1150 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1150 <= regs_1149; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1151 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1151 <= regs_1150; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1152 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1152 <= regs_1151; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1153 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1153 <= regs_1152; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1154 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1154 <= regs_1153; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1155 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1155 <= regs_1154; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1156 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1156 <= regs_1155; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1157 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1157 <= regs_1156; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1158 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1158 <= regs_1157; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1159 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1159 <= regs_1158; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1160 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1160 <= regs_1159; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1161 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1161 <= regs_1160; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1162 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1162 <= regs_1161; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1163 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1163 <= regs_1162; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1164 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1164 <= regs_1163; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1165 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1165 <= regs_1164; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1166 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1166 <= regs_1165; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1167 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1167 <= regs_1166; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1168 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1168 <= regs_1167; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1169 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1169 <= regs_1168; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1170 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1170 <= regs_1169; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1171 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1171 <= regs_1170; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1172 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1172 <= regs_1171; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1173 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1173 <= regs_1172; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1174 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1174 <= regs_1173; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1175 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1175 <= regs_1174; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1176 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1176 <= regs_1175; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1177 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1177 <= regs_1176; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1178 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1178 <= regs_1177; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1179 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1179 <= regs_1178; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1180 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1180 <= regs_1179; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1181 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1181 <= regs_1180; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1182 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1182 <= regs_1181; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1183 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1183 <= regs_1182; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1184 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1184 <= regs_1183; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1185 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1185 <= regs_1184; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1186 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1186 <= regs_1185; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1187 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1187 <= regs_1186; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1188 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1188 <= regs_1187; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1189 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1189 <= regs_1188; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1190 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1190 <= regs_1189; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1191 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1191 <= regs_1190; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1192 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1192 <= regs_1191; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1193 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1193 <= regs_1192; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1194 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1194 <= regs_1193; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1195 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1195 <= regs_1194; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1196 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1196 <= regs_1195; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1197 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1197 <= regs_1196; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1198 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1198 <= regs_1197; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1199 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1199 <= regs_1198; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1200 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1200 <= regs_1199; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1201 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1201 <= regs_1200; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1202 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1202 <= regs_1201; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1203 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1203 <= regs_1202; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1204 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1204 <= regs_1203; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1205 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1205 <= regs_1204; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1206 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1206 <= regs_1205; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1207 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1207 <= regs_1206; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1208 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1208 <= regs_1207; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1209 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1209 <= regs_1208; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1210 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1210 <= regs_1209; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1211 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1211 <= regs_1210; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1212 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1212 <= regs_1211; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1213 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1213 <= regs_1212; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1214 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1214 <= regs_1213; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1215 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1215 <= regs_1214; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1216 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1216 <= regs_1215; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1217 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1217 <= regs_1216; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1218 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1218 <= regs_1217; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1219 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1219 <= regs_1218; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1220 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1220 <= regs_1219; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1221 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1221 <= regs_1220; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1222 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1222 <= regs_1221; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1223 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1223 <= regs_1222; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1224 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1224 <= regs_1223; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1225 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1225 <= regs_1224; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1226 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1226 <= regs_1225; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1227 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1227 <= regs_1226; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1228 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1228 <= regs_1227; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1229 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1229 <= regs_1228; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1230 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1230 <= regs_1229; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1231 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1231 <= regs_1230; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1232 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1232 <= regs_1231; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1233 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1233 <= regs_1232; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1234 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1234 <= regs_1233; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1235 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1235 <= regs_1234; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1236 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1236 <= regs_1235; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1237 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1237 <= regs_1236; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1238 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1238 <= regs_1237; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1239 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1239 <= regs_1238; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1240 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1240 <= regs_1239; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1241 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1241 <= regs_1240; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1242 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1242 <= regs_1241; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1243 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1243 <= regs_1242; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1244 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1244 <= regs_1243; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1245 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1245 <= regs_1244; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1246 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1246 <= regs_1245; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1247 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1247 <= regs_1246; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1248 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1248 <= regs_1247; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1249 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1249 <= regs_1248; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1250 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1250 <= regs_1249; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1251 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1251 <= regs_1250; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1252 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1252 <= regs_1251; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1253 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1253 <= regs_1252; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1254 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1254 <= regs_1253; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1255 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1255 <= regs_1254; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1256 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1256 <= regs_1255; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1257 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1257 <= regs_1256; // @[FloatingPointDesigns.scala 2277:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2274:23]
      regs_1258 <= 32'h0; // @[FloatingPointDesigns.scala 2274:23]
    end else begin
      regs_1258 <= regs_1257; // @[FloatingPointDesigns.scala 2277:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  regs_64 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  regs_65 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  regs_66 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  regs_67 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  regs_68 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  regs_69 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  regs_70 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  regs_71 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  regs_72 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  regs_73 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  regs_74 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  regs_75 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  regs_76 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  regs_77 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  regs_78 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  regs_79 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  regs_80 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  regs_81 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  regs_82 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  regs_83 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  regs_84 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  regs_85 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  regs_86 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  regs_87 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  regs_88 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  regs_89 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  regs_90 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  regs_91 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  regs_92 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  regs_93 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  regs_94 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  regs_95 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  regs_96 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  regs_97 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  regs_98 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  regs_99 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  regs_100 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  regs_101 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  regs_102 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  regs_103 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  regs_104 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  regs_105 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  regs_106 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  regs_107 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  regs_108 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  regs_109 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  regs_110 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  regs_111 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  regs_112 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  regs_113 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  regs_114 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  regs_115 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  regs_116 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  regs_117 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  regs_118 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  regs_119 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  regs_120 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  regs_121 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  regs_122 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  regs_123 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  regs_124 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  regs_125 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  regs_126 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  regs_127 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  regs_128 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  regs_129 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  regs_130 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  regs_131 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  regs_132 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  regs_133 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  regs_134 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  regs_135 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  regs_136 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  regs_137 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  regs_138 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  regs_139 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  regs_140 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  regs_141 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  regs_142 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  regs_143 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  regs_144 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  regs_145 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  regs_146 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  regs_147 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  regs_148 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  regs_149 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  regs_150 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  regs_151 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  regs_152 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  regs_153 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  regs_154 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  regs_155 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  regs_156 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  regs_157 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  regs_158 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  regs_159 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  regs_160 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  regs_161 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  regs_162 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  regs_163 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  regs_164 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  regs_165 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  regs_166 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  regs_167 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  regs_168 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  regs_169 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  regs_170 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  regs_171 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  regs_172 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  regs_173 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  regs_174 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  regs_175 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  regs_176 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  regs_177 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  regs_178 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  regs_179 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  regs_180 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  regs_181 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  regs_182 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  regs_183 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  regs_184 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  regs_185 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  regs_186 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  regs_187 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  regs_188 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  regs_189 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  regs_190 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  regs_191 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  regs_192 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  regs_193 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  regs_194 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  regs_195 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  regs_196 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  regs_197 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  regs_198 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  regs_199 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  regs_200 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  regs_201 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  regs_202 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  regs_203 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  regs_204 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  regs_205 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  regs_206 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  regs_207 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  regs_208 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  regs_209 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  regs_210 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  regs_211 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  regs_212 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  regs_213 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  regs_214 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  regs_215 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  regs_216 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  regs_217 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  regs_218 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  regs_219 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  regs_220 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  regs_221 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  regs_222 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  regs_223 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  regs_224 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  regs_225 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  regs_226 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  regs_227 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  regs_228 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  regs_229 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  regs_230 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  regs_231 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  regs_232 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  regs_233 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  regs_234 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  regs_235 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  regs_236 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  regs_237 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  regs_238 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  regs_239 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  regs_240 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  regs_241 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  regs_242 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  regs_243 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  regs_244 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  regs_245 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  regs_246 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  regs_247 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  regs_248 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  regs_249 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  regs_250 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  regs_251 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  regs_252 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  regs_253 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  regs_254 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  regs_255 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  regs_256 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  regs_257 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  regs_258 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  regs_259 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  regs_260 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  regs_261 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  regs_262 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  regs_263 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  regs_264 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  regs_265 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  regs_266 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  regs_267 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  regs_268 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  regs_269 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  regs_270 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  regs_271 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  regs_272 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  regs_273 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  regs_274 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  regs_275 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  regs_276 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  regs_277 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  regs_278 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  regs_279 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  regs_280 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  regs_281 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  regs_282 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  regs_283 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  regs_284 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  regs_285 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  regs_286 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  regs_287 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  regs_288 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  regs_289 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  regs_290 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  regs_291 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  regs_292 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  regs_293 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  regs_294 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  regs_295 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  regs_296 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  regs_297 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  regs_298 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  regs_299 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  regs_300 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  regs_301 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  regs_302 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  regs_303 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  regs_304 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  regs_305 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  regs_306 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  regs_307 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  regs_308 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  regs_309 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  regs_310 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  regs_311 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  regs_312 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  regs_313 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  regs_314 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  regs_315 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  regs_316 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  regs_317 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  regs_318 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  regs_319 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  regs_320 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  regs_321 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  regs_322 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  regs_323 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  regs_324 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  regs_325 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  regs_326 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  regs_327 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  regs_328 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  regs_329 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  regs_330 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  regs_331 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  regs_332 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  regs_333 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  regs_334 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  regs_335 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  regs_336 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  regs_337 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  regs_338 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  regs_339 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  regs_340 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  regs_341 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  regs_342 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  regs_343 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  regs_344 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  regs_345 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  regs_346 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  regs_347 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  regs_348 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  regs_349 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  regs_350 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  regs_351 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  regs_352 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  regs_353 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  regs_354 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  regs_355 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  regs_356 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  regs_357 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  regs_358 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  regs_359 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  regs_360 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  regs_361 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  regs_362 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  regs_363 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  regs_364 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  regs_365 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  regs_366 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  regs_367 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  regs_368 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  regs_369 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  regs_370 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  regs_371 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  regs_372 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  regs_373 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  regs_374 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  regs_375 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  regs_376 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  regs_377 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  regs_378 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  regs_379 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  regs_380 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  regs_381 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  regs_382 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  regs_383 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  regs_384 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  regs_385 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  regs_386 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  regs_387 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  regs_388 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  regs_389 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  regs_390 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  regs_391 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  regs_392 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  regs_393 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  regs_394 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  regs_395 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  regs_396 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  regs_397 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  regs_398 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  regs_399 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  regs_400 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  regs_401 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  regs_402 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  regs_403 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  regs_404 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  regs_405 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  regs_406 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  regs_407 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  regs_408 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  regs_409 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  regs_410 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  regs_411 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  regs_412 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  regs_413 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  regs_414 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  regs_415 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  regs_416 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  regs_417 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  regs_418 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  regs_419 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  regs_420 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  regs_421 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  regs_422 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  regs_423 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  regs_424 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  regs_425 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  regs_426 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  regs_427 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  regs_428 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  regs_429 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  regs_430 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  regs_431 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  regs_432 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  regs_433 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  regs_434 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  regs_435 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  regs_436 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  regs_437 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  regs_438 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  regs_439 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  regs_440 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  regs_441 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  regs_442 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  regs_443 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  regs_444 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  regs_445 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  regs_446 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  regs_447 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  regs_448 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  regs_449 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  regs_450 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  regs_451 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  regs_452 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  regs_453 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  regs_454 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  regs_455 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  regs_456 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  regs_457 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  regs_458 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  regs_459 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  regs_460 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  regs_461 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  regs_462 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  regs_463 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  regs_464 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  regs_465 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  regs_466 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  regs_467 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  regs_468 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  regs_469 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  regs_470 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  regs_471 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  regs_472 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  regs_473 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  regs_474 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  regs_475 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  regs_476 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  regs_477 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  regs_478 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  regs_479 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  regs_480 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  regs_481 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  regs_482 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  regs_483 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  regs_484 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  regs_485 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  regs_486 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  regs_487 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  regs_488 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  regs_489 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  regs_490 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  regs_491 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  regs_492 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  regs_493 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  regs_494 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  regs_495 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  regs_496 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  regs_497 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  regs_498 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  regs_499 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  regs_500 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  regs_501 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  regs_502 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  regs_503 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  regs_504 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  regs_505 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  regs_506 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  regs_507 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  regs_508 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  regs_509 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  regs_510 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  regs_511 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  regs_512 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  regs_513 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  regs_514 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  regs_515 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  regs_516 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  regs_517 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  regs_518 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  regs_519 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  regs_520 = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  regs_521 = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  regs_522 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  regs_523 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  regs_524 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  regs_525 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  regs_526 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  regs_527 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  regs_528 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  regs_529 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  regs_530 = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  regs_531 = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  regs_532 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  regs_533 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  regs_534 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  regs_535 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  regs_536 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  regs_537 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  regs_538 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  regs_539 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  regs_540 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  regs_541 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  regs_542 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  regs_543 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  regs_544 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  regs_545 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  regs_546 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  regs_547 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  regs_548 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  regs_549 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  regs_550 = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  regs_551 = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  regs_552 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  regs_553 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  regs_554 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  regs_555 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  regs_556 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  regs_557 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  regs_558 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  regs_559 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  regs_560 = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  regs_561 = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  regs_562 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  regs_563 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  regs_564 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  regs_565 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  regs_566 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  regs_567 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  regs_568 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  regs_569 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  regs_570 = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  regs_571 = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  regs_572 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  regs_573 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  regs_574 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  regs_575 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  regs_576 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  regs_577 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  regs_578 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  regs_579 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  regs_580 = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  regs_581 = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  regs_582 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  regs_583 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  regs_584 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  regs_585 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  regs_586 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  regs_587 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  regs_588 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  regs_589 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  regs_590 = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  regs_591 = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  regs_592 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  regs_593 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  regs_594 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  regs_595 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  regs_596 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  regs_597 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  regs_598 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  regs_599 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  regs_600 = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  regs_601 = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  regs_602 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  regs_603 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  regs_604 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  regs_605 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  regs_606 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  regs_607 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  regs_608 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  regs_609 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  regs_610 = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  regs_611 = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  regs_612 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  regs_613 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  regs_614 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  regs_615 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  regs_616 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  regs_617 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  regs_618 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  regs_619 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  regs_620 = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  regs_621 = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  regs_622 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  regs_623 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  regs_624 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  regs_625 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  regs_626 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  regs_627 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  regs_628 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  regs_629 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  regs_630 = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  regs_631 = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  regs_632 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  regs_633 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  regs_634 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  regs_635 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  regs_636 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  regs_637 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  regs_638 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  regs_639 = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  regs_640 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  regs_641 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  regs_642 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  regs_643 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  regs_644 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  regs_645 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  regs_646 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  regs_647 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  regs_648 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  regs_649 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  regs_650 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  regs_651 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  regs_652 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  regs_653 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  regs_654 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  regs_655 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  regs_656 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  regs_657 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  regs_658 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  regs_659 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  regs_660 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  regs_661 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  regs_662 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  regs_663 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  regs_664 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  regs_665 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  regs_666 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  regs_667 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  regs_668 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  regs_669 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  regs_670 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  regs_671 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  regs_672 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  regs_673 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  regs_674 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  regs_675 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  regs_676 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  regs_677 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  regs_678 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  regs_679 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  regs_680 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  regs_681 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  regs_682 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  regs_683 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  regs_684 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  regs_685 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  regs_686 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  regs_687 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  regs_688 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  regs_689 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  regs_690 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  regs_691 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  regs_692 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  regs_693 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  regs_694 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  regs_695 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  regs_696 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  regs_697 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  regs_698 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  regs_699 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  regs_700 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  regs_701 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  regs_702 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  regs_703 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  regs_704 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  regs_705 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  regs_706 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  regs_707 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  regs_708 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  regs_709 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  regs_710 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  regs_711 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  regs_712 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  regs_713 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  regs_714 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  regs_715 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  regs_716 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  regs_717 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  regs_718 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  regs_719 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  regs_720 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  regs_721 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  regs_722 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  regs_723 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  regs_724 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  regs_725 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  regs_726 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  regs_727 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  regs_728 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  regs_729 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  regs_730 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  regs_731 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  regs_732 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  regs_733 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  regs_734 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  regs_735 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  regs_736 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  regs_737 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  regs_738 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  regs_739 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  regs_740 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  regs_741 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  regs_742 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  regs_743 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  regs_744 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  regs_745 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  regs_746 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  regs_747 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  regs_748 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  regs_749 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  regs_750 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  regs_751 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  regs_752 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  regs_753 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  regs_754 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  regs_755 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  regs_756 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  regs_757 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  regs_758 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  regs_759 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  regs_760 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  regs_761 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  regs_762 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  regs_763 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  regs_764 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  regs_765 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  regs_766 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  regs_767 = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  regs_768 = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  regs_769 = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  regs_770 = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  regs_771 = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  regs_772 = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  regs_773 = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  regs_774 = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  regs_775 = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  regs_776 = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  regs_777 = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  regs_778 = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  regs_779 = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  regs_780 = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  regs_781 = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  regs_782 = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  regs_783 = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  regs_784 = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  regs_785 = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  regs_786 = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  regs_787 = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  regs_788 = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  regs_789 = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  regs_790 = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  regs_791 = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  regs_792 = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  regs_793 = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  regs_794 = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  regs_795 = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  regs_796 = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  regs_797 = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  regs_798 = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  regs_799 = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  regs_800 = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  regs_801 = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  regs_802 = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  regs_803 = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  regs_804 = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  regs_805 = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  regs_806 = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  regs_807 = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  regs_808 = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  regs_809 = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  regs_810 = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  regs_811 = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  regs_812 = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  regs_813 = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  regs_814 = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  regs_815 = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  regs_816 = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  regs_817 = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  regs_818 = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  regs_819 = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  regs_820 = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  regs_821 = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  regs_822 = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  regs_823 = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  regs_824 = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  regs_825 = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  regs_826 = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  regs_827 = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  regs_828 = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  regs_829 = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  regs_830 = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  regs_831 = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  regs_832 = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  regs_833 = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  regs_834 = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  regs_835 = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  regs_836 = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  regs_837 = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  regs_838 = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  regs_839 = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  regs_840 = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  regs_841 = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  regs_842 = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  regs_843 = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  regs_844 = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  regs_845 = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  regs_846 = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  regs_847 = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  regs_848 = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  regs_849 = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  regs_850 = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  regs_851 = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  regs_852 = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  regs_853 = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  regs_854 = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  regs_855 = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  regs_856 = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  regs_857 = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  regs_858 = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  regs_859 = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  regs_860 = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  regs_861 = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  regs_862 = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  regs_863 = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  regs_864 = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  regs_865 = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  regs_866 = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  regs_867 = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  regs_868 = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  regs_869 = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  regs_870 = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  regs_871 = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  regs_872 = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  regs_873 = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  regs_874 = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  regs_875 = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  regs_876 = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  regs_877 = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  regs_878 = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  regs_879 = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  regs_880 = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  regs_881 = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  regs_882 = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  regs_883 = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  regs_884 = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  regs_885 = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  regs_886 = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  regs_887 = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  regs_888 = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  regs_889 = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  regs_890 = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  regs_891 = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  regs_892 = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  regs_893 = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  regs_894 = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  regs_895 = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  regs_896 = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  regs_897 = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  regs_898 = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  regs_899 = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  regs_900 = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  regs_901 = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  regs_902 = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  regs_903 = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  regs_904 = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  regs_905 = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  regs_906 = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  regs_907 = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  regs_908 = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  regs_909 = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  regs_910 = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  regs_911 = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  regs_912 = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  regs_913 = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  regs_914 = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  regs_915 = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  regs_916 = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  regs_917 = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  regs_918 = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  regs_919 = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  regs_920 = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  regs_921 = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  regs_922 = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  regs_923 = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  regs_924 = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  regs_925 = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  regs_926 = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  regs_927 = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  regs_928 = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  regs_929 = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  regs_930 = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  regs_931 = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  regs_932 = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  regs_933 = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  regs_934 = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  regs_935 = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  regs_936 = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  regs_937 = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  regs_938 = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  regs_939 = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  regs_940 = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  regs_941 = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  regs_942 = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  regs_943 = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  regs_944 = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  regs_945 = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  regs_946 = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  regs_947 = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  regs_948 = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  regs_949 = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  regs_950 = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  regs_951 = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  regs_952 = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  regs_953 = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  regs_954 = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  regs_955 = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  regs_956 = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  regs_957 = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  regs_958 = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  regs_959 = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  regs_960 = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  regs_961 = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  regs_962 = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  regs_963 = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  regs_964 = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  regs_965 = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  regs_966 = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  regs_967 = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  regs_968 = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  regs_969 = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  regs_970 = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  regs_971 = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  regs_972 = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  regs_973 = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  regs_974 = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  regs_975 = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  regs_976 = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  regs_977 = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  regs_978 = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  regs_979 = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  regs_980 = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  regs_981 = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  regs_982 = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  regs_983 = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  regs_984 = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  regs_985 = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  regs_986 = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  regs_987 = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  regs_988 = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  regs_989 = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  regs_990 = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  regs_991 = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  regs_992 = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  regs_993 = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  regs_994 = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  regs_995 = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  regs_996 = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  regs_997 = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  regs_998 = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  regs_999 = _RAND_999[31:0];
  _RAND_1000 = {1{`RANDOM}};
  regs_1000 = _RAND_1000[31:0];
  _RAND_1001 = {1{`RANDOM}};
  regs_1001 = _RAND_1001[31:0];
  _RAND_1002 = {1{`RANDOM}};
  regs_1002 = _RAND_1002[31:0];
  _RAND_1003 = {1{`RANDOM}};
  regs_1003 = _RAND_1003[31:0];
  _RAND_1004 = {1{`RANDOM}};
  regs_1004 = _RAND_1004[31:0];
  _RAND_1005 = {1{`RANDOM}};
  regs_1005 = _RAND_1005[31:0];
  _RAND_1006 = {1{`RANDOM}};
  regs_1006 = _RAND_1006[31:0];
  _RAND_1007 = {1{`RANDOM}};
  regs_1007 = _RAND_1007[31:0];
  _RAND_1008 = {1{`RANDOM}};
  regs_1008 = _RAND_1008[31:0];
  _RAND_1009 = {1{`RANDOM}};
  regs_1009 = _RAND_1009[31:0];
  _RAND_1010 = {1{`RANDOM}};
  regs_1010 = _RAND_1010[31:0];
  _RAND_1011 = {1{`RANDOM}};
  regs_1011 = _RAND_1011[31:0];
  _RAND_1012 = {1{`RANDOM}};
  regs_1012 = _RAND_1012[31:0];
  _RAND_1013 = {1{`RANDOM}};
  regs_1013 = _RAND_1013[31:0];
  _RAND_1014 = {1{`RANDOM}};
  regs_1014 = _RAND_1014[31:0];
  _RAND_1015 = {1{`RANDOM}};
  regs_1015 = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  regs_1016 = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  regs_1017 = _RAND_1017[31:0];
  _RAND_1018 = {1{`RANDOM}};
  regs_1018 = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  regs_1019 = _RAND_1019[31:0];
  _RAND_1020 = {1{`RANDOM}};
  regs_1020 = _RAND_1020[31:0];
  _RAND_1021 = {1{`RANDOM}};
  regs_1021 = _RAND_1021[31:0];
  _RAND_1022 = {1{`RANDOM}};
  regs_1022 = _RAND_1022[31:0];
  _RAND_1023 = {1{`RANDOM}};
  regs_1023 = _RAND_1023[31:0];
  _RAND_1024 = {1{`RANDOM}};
  regs_1024 = _RAND_1024[31:0];
  _RAND_1025 = {1{`RANDOM}};
  regs_1025 = _RAND_1025[31:0];
  _RAND_1026 = {1{`RANDOM}};
  regs_1026 = _RAND_1026[31:0];
  _RAND_1027 = {1{`RANDOM}};
  regs_1027 = _RAND_1027[31:0];
  _RAND_1028 = {1{`RANDOM}};
  regs_1028 = _RAND_1028[31:0];
  _RAND_1029 = {1{`RANDOM}};
  regs_1029 = _RAND_1029[31:0];
  _RAND_1030 = {1{`RANDOM}};
  regs_1030 = _RAND_1030[31:0];
  _RAND_1031 = {1{`RANDOM}};
  regs_1031 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  regs_1032 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  regs_1033 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  regs_1034 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  regs_1035 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  regs_1036 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  regs_1037 = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  regs_1038 = _RAND_1038[31:0];
  _RAND_1039 = {1{`RANDOM}};
  regs_1039 = _RAND_1039[31:0];
  _RAND_1040 = {1{`RANDOM}};
  regs_1040 = _RAND_1040[31:0];
  _RAND_1041 = {1{`RANDOM}};
  regs_1041 = _RAND_1041[31:0];
  _RAND_1042 = {1{`RANDOM}};
  regs_1042 = _RAND_1042[31:0];
  _RAND_1043 = {1{`RANDOM}};
  regs_1043 = _RAND_1043[31:0];
  _RAND_1044 = {1{`RANDOM}};
  regs_1044 = _RAND_1044[31:0];
  _RAND_1045 = {1{`RANDOM}};
  regs_1045 = _RAND_1045[31:0];
  _RAND_1046 = {1{`RANDOM}};
  regs_1046 = _RAND_1046[31:0];
  _RAND_1047 = {1{`RANDOM}};
  regs_1047 = _RAND_1047[31:0];
  _RAND_1048 = {1{`RANDOM}};
  regs_1048 = _RAND_1048[31:0];
  _RAND_1049 = {1{`RANDOM}};
  regs_1049 = _RAND_1049[31:0];
  _RAND_1050 = {1{`RANDOM}};
  regs_1050 = _RAND_1050[31:0];
  _RAND_1051 = {1{`RANDOM}};
  regs_1051 = _RAND_1051[31:0];
  _RAND_1052 = {1{`RANDOM}};
  regs_1052 = _RAND_1052[31:0];
  _RAND_1053 = {1{`RANDOM}};
  regs_1053 = _RAND_1053[31:0];
  _RAND_1054 = {1{`RANDOM}};
  regs_1054 = _RAND_1054[31:0];
  _RAND_1055 = {1{`RANDOM}};
  regs_1055 = _RAND_1055[31:0];
  _RAND_1056 = {1{`RANDOM}};
  regs_1056 = _RAND_1056[31:0];
  _RAND_1057 = {1{`RANDOM}};
  regs_1057 = _RAND_1057[31:0];
  _RAND_1058 = {1{`RANDOM}};
  regs_1058 = _RAND_1058[31:0];
  _RAND_1059 = {1{`RANDOM}};
  regs_1059 = _RAND_1059[31:0];
  _RAND_1060 = {1{`RANDOM}};
  regs_1060 = _RAND_1060[31:0];
  _RAND_1061 = {1{`RANDOM}};
  regs_1061 = _RAND_1061[31:0];
  _RAND_1062 = {1{`RANDOM}};
  regs_1062 = _RAND_1062[31:0];
  _RAND_1063 = {1{`RANDOM}};
  regs_1063 = _RAND_1063[31:0];
  _RAND_1064 = {1{`RANDOM}};
  regs_1064 = _RAND_1064[31:0];
  _RAND_1065 = {1{`RANDOM}};
  regs_1065 = _RAND_1065[31:0];
  _RAND_1066 = {1{`RANDOM}};
  regs_1066 = _RAND_1066[31:0];
  _RAND_1067 = {1{`RANDOM}};
  regs_1067 = _RAND_1067[31:0];
  _RAND_1068 = {1{`RANDOM}};
  regs_1068 = _RAND_1068[31:0];
  _RAND_1069 = {1{`RANDOM}};
  regs_1069 = _RAND_1069[31:0];
  _RAND_1070 = {1{`RANDOM}};
  regs_1070 = _RAND_1070[31:0];
  _RAND_1071 = {1{`RANDOM}};
  regs_1071 = _RAND_1071[31:0];
  _RAND_1072 = {1{`RANDOM}};
  regs_1072 = _RAND_1072[31:0];
  _RAND_1073 = {1{`RANDOM}};
  regs_1073 = _RAND_1073[31:0];
  _RAND_1074 = {1{`RANDOM}};
  regs_1074 = _RAND_1074[31:0];
  _RAND_1075 = {1{`RANDOM}};
  regs_1075 = _RAND_1075[31:0];
  _RAND_1076 = {1{`RANDOM}};
  regs_1076 = _RAND_1076[31:0];
  _RAND_1077 = {1{`RANDOM}};
  regs_1077 = _RAND_1077[31:0];
  _RAND_1078 = {1{`RANDOM}};
  regs_1078 = _RAND_1078[31:0];
  _RAND_1079 = {1{`RANDOM}};
  regs_1079 = _RAND_1079[31:0];
  _RAND_1080 = {1{`RANDOM}};
  regs_1080 = _RAND_1080[31:0];
  _RAND_1081 = {1{`RANDOM}};
  regs_1081 = _RAND_1081[31:0];
  _RAND_1082 = {1{`RANDOM}};
  regs_1082 = _RAND_1082[31:0];
  _RAND_1083 = {1{`RANDOM}};
  regs_1083 = _RAND_1083[31:0];
  _RAND_1084 = {1{`RANDOM}};
  regs_1084 = _RAND_1084[31:0];
  _RAND_1085 = {1{`RANDOM}};
  regs_1085 = _RAND_1085[31:0];
  _RAND_1086 = {1{`RANDOM}};
  regs_1086 = _RAND_1086[31:0];
  _RAND_1087 = {1{`RANDOM}};
  regs_1087 = _RAND_1087[31:0];
  _RAND_1088 = {1{`RANDOM}};
  regs_1088 = _RAND_1088[31:0];
  _RAND_1089 = {1{`RANDOM}};
  regs_1089 = _RAND_1089[31:0];
  _RAND_1090 = {1{`RANDOM}};
  regs_1090 = _RAND_1090[31:0];
  _RAND_1091 = {1{`RANDOM}};
  regs_1091 = _RAND_1091[31:0];
  _RAND_1092 = {1{`RANDOM}};
  regs_1092 = _RAND_1092[31:0];
  _RAND_1093 = {1{`RANDOM}};
  regs_1093 = _RAND_1093[31:0];
  _RAND_1094 = {1{`RANDOM}};
  regs_1094 = _RAND_1094[31:0];
  _RAND_1095 = {1{`RANDOM}};
  regs_1095 = _RAND_1095[31:0];
  _RAND_1096 = {1{`RANDOM}};
  regs_1096 = _RAND_1096[31:0];
  _RAND_1097 = {1{`RANDOM}};
  regs_1097 = _RAND_1097[31:0];
  _RAND_1098 = {1{`RANDOM}};
  regs_1098 = _RAND_1098[31:0];
  _RAND_1099 = {1{`RANDOM}};
  regs_1099 = _RAND_1099[31:0];
  _RAND_1100 = {1{`RANDOM}};
  regs_1100 = _RAND_1100[31:0];
  _RAND_1101 = {1{`RANDOM}};
  regs_1101 = _RAND_1101[31:0];
  _RAND_1102 = {1{`RANDOM}};
  regs_1102 = _RAND_1102[31:0];
  _RAND_1103 = {1{`RANDOM}};
  regs_1103 = _RAND_1103[31:0];
  _RAND_1104 = {1{`RANDOM}};
  regs_1104 = _RAND_1104[31:0];
  _RAND_1105 = {1{`RANDOM}};
  regs_1105 = _RAND_1105[31:0];
  _RAND_1106 = {1{`RANDOM}};
  regs_1106 = _RAND_1106[31:0];
  _RAND_1107 = {1{`RANDOM}};
  regs_1107 = _RAND_1107[31:0];
  _RAND_1108 = {1{`RANDOM}};
  regs_1108 = _RAND_1108[31:0];
  _RAND_1109 = {1{`RANDOM}};
  regs_1109 = _RAND_1109[31:0];
  _RAND_1110 = {1{`RANDOM}};
  regs_1110 = _RAND_1110[31:0];
  _RAND_1111 = {1{`RANDOM}};
  regs_1111 = _RAND_1111[31:0];
  _RAND_1112 = {1{`RANDOM}};
  regs_1112 = _RAND_1112[31:0];
  _RAND_1113 = {1{`RANDOM}};
  regs_1113 = _RAND_1113[31:0];
  _RAND_1114 = {1{`RANDOM}};
  regs_1114 = _RAND_1114[31:0];
  _RAND_1115 = {1{`RANDOM}};
  regs_1115 = _RAND_1115[31:0];
  _RAND_1116 = {1{`RANDOM}};
  regs_1116 = _RAND_1116[31:0];
  _RAND_1117 = {1{`RANDOM}};
  regs_1117 = _RAND_1117[31:0];
  _RAND_1118 = {1{`RANDOM}};
  regs_1118 = _RAND_1118[31:0];
  _RAND_1119 = {1{`RANDOM}};
  regs_1119 = _RAND_1119[31:0];
  _RAND_1120 = {1{`RANDOM}};
  regs_1120 = _RAND_1120[31:0];
  _RAND_1121 = {1{`RANDOM}};
  regs_1121 = _RAND_1121[31:0];
  _RAND_1122 = {1{`RANDOM}};
  regs_1122 = _RAND_1122[31:0];
  _RAND_1123 = {1{`RANDOM}};
  regs_1123 = _RAND_1123[31:0];
  _RAND_1124 = {1{`RANDOM}};
  regs_1124 = _RAND_1124[31:0];
  _RAND_1125 = {1{`RANDOM}};
  regs_1125 = _RAND_1125[31:0];
  _RAND_1126 = {1{`RANDOM}};
  regs_1126 = _RAND_1126[31:0];
  _RAND_1127 = {1{`RANDOM}};
  regs_1127 = _RAND_1127[31:0];
  _RAND_1128 = {1{`RANDOM}};
  regs_1128 = _RAND_1128[31:0];
  _RAND_1129 = {1{`RANDOM}};
  regs_1129 = _RAND_1129[31:0];
  _RAND_1130 = {1{`RANDOM}};
  regs_1130 = _RAND_1130[31:0];
  _RAND_1131 = {1{`RANDOM}};
  regs_1131 = _RAND_1131[31:0];
  _RAND_1132 = {1{`RANDOM}};
  regs_1132 = _RAND_1132[31:0];
  _RAND_1133 = {1{`RANDOM}};
  regs_1133 = _RAND_1133[31:0];
  _RAND_1134 = {1{`RANDOM}};
  regs_1134 = _RAND_1134[31:0];
  _RAND_1135 = {1{`RANDOM}};
  regs_1135 = _RAND_1135[31:0];
  _RAND_1136 = {1{`RANDOM}};
  regs_1136 = _RAND_1136[31:0];
  _RAND_1137 = {1{`RANDOM}};
  regs_1137 = _RAND_1137[31:0];
  _RAND_1138 = {1{`RANDOM}};
  regs_1138 = _RAND_1138[31:0];
  _RAND_1139 = {1{`RANDOM}};
  regs_1139 = _RAND_1139[31:0];
  _RAND_1140 = {1{`RANDOM}};
  regs_1140 = _RAND_1140[31:0];
  _RAND_1141 = {1{`RANDOM}};
  regs_1141 = _RAND_1141[31:0];
  _RAND_1142 = {1{`RANDOM}};
  regs_1142 = _RAND_1142[31:0];
  _RAND_1143 = {1{`RANDOM}};
  regs_1143 = _RAND_1143[31:0];
  _RAND_1144 = {1{`RANDOM}};
  regs_1144 = _RAND_1144[31:0];
  _RAND_1145 = {1{`RANDOM}};
  regs_1145 = _RAND_1145[31:0];
  _RAND_1146 = {1{`RANDOM}};
  regs_1146 = _RAND_1146[31:0];
  _RAND_1147 = {1{`RANDOM}};
  regs_1147 = _RAND_1147[31:0];
  _RAND_1148 = {1{`RANDOM}};
  regs_1148 = _RAND_1148[31:0];
  _RAND_1149 = {1{`RANDOM}};
  regs_1149 = _RAND_1149[31:0];
  _RAND_1150 = {1{`RANDOM}};
  regs_1150 = _RAND_1150[31:0];
  _RAND_1151 = {1{`RANDOM}};
  regs_1151 = _RAND_1151[31:0];
  _RAND_1152 = {1{`RANDOM}};
  regs_1152 = _RAND_1152[31:0];
  _RAND_1153 = {1{`RANDOM}};
  regs_1153 = _RAND_1153[31:0];
  _RAND_1154 = {1{`RANDOM}};
  regs_1154 = _RAND_1154[31:0];
  _RAND_1155 = {1{`RANDOM}};
  regs_1155 = _RAND_1155[31:0];
  _RAND_1156 = {1{`RANDOM}};
  regs_1156 = _RAND_1156[31:0];
  _RAND_1157 = {1{`RANDOM}};
  regs_1157 = _RAND_1157[31:0];
  _RAND_1158 = {1{`RANDOM}};
  regs_1158 = _RAND_1158[31:0];
  _RAND_1159 = {1{`RANDOM}};
  regs_1159 = _RAND_1159[31:0];
  _RAND_1160 = {1{`RANDOM}};
  regs_1160 = _RAND_1160[31:0];
  _RAND_1161 = {1{`RANDOM}};
  regs_1161 = _RAND_1161[31:0];
  _RAND_1162 = {1{`RANDOM}};
  regs_1162 = _RAND_1162[31:0];
  _RAND_1163 = {1{`RANDOM}};
  regs_1163 = _RAND_1163[31:0];
  _RAND_1164 = {1{`RANDOM}};
  regs_1164 = _RAND_1164[31:0];
  _RAND_1165 = {1{`RANDOM}};
  regs_1165 = _RAND_1165[31:0];
  _RAND_1166 = {1{`RANDOM}};
  regs_1166 = _RAND_1166[31:0];
  _RAND_1167 = {1{`RANDOM}};
  regs_1167 = _RAND_1167[31:0];
  _RAND_1168 = {1{`RANDOM}};
  regs_1168 = _RAND_1168[31:0];
  _RAND_1169 = {1{`RANDOM}};
  regs_1169 = _RAND_1169[31:0];
  _RAND_1170 = {1{`RANDOM}};
  regs_1170 = _RAND_1170[31:0];
  _RAND_1171 = {1{`RANDOM}};
  regs_1171 = _RAND_1171[31:0];
  _RAND_1172 = {1{`RANDOM}};
  regs_1172 = _RAND_1172[31:0];
  _RAND_1173 = {1{`RANDOM}};
  regs_1173 = _RAND_1173[31:0];
  _RAND_1174 = {1{`RANDOM}};
  regs_1174 = _RAND_1174[31:0];
  _RAND_1175 = {1{`RANDOM}};
  regs_1175 = _RAND_1175[31:0];
  _RAND_1176 = {1{`RANDOM}};
  regs_1176 = _RAND_1176[31:0];
  _RAND_1177 = {1{`RANDOM}};
  regs_1177 = _RAND_1177[31:0];
  _RAND_1178 = {1{`RANDOM}};
  regs_1178 = _RAND_1178[31:0];
  _RAND_1179 = {1{`RANDOM}};
  regs_1179 = _RAND_1179[31:0];
  _RAND_1180 = {1{`RANDOM}};
  regs_1180 = _RAND_1180[31:0];
  _RAND_1181 = {1{`RANDOM}};
  regs_1181 = _RAND_1181[31:0];
  _RAND_1182 = {1{`RANDOM}};
  regs_1182 = _RAND_1182[31:0];
  _RAND_1183 = {1{`RANDOM}};
  regs_1183 = _RAND_1183[31:0];
  _RAND_1184 = {1{`RANDOM}};
  regs_1184 = _RAND_1184[31:0];
  _RAND_1185 = {1{`RANDOM}};
  regs_1185 = _RAND_1185[31:0];
  _RAND_1186 = {1{`RANDOM}};
  regs_1186 = _RAND_1186[31:0];
  _RAND_1187 = {1{`RANDOM}};
  regs_1187 = _RAND_1187[31:0];
  _RAND_1188 = {1{`RANDOM}};
  regs_1188 = _RAND_1188[31:0];
  _RAND_1189 = {1{`RANDOM}};
  regs_1189 = _RAND_1189[31:0];
  _RAND_1190 = {1{`RANDOM}};
  regs_1190 = _RAND_1190[31:0];
  _RAND_1191 = {1{`RANDOM}};
  regs_1191 = _RAND_1191[31:0];
  _RAND_1192 = {1{`RANDOM}};
  regs_1192 = _RAND_1192[31:0];
  _RAND_1193 = {1{`RANDOM}};
  regs_1193 = _RAND_1193[31:0];
  _RAND_1194 = {1{`RANDOM}};
  regs_1194 = _RAND_1194[31:0];
  _RAND_1195 = {1{`RANDOM}};
  regs_1195 = _RAND_1195[31:0];
  _RAND_1196 = {1{`RANDOM}};
  regs_1196 = _RAND_1196[31:0];
  _RAND_1197 = {1{`RANDOM}};
  regs_1197 = _RAND_1197[31:0];
  _RAND_1198 = {1{`RANDOM}};
  regs_1198 = _RAND_1198[31:0];
  _RAND_1199 = {1{`RANDOM}};
  regs_1199 = _RAND_1199[31:0];
  _RAND_1200 = {1{`RANDOM}};
  regs_1200 = _RAND_1200[31:0];
  _RAND_1201 = {1{`RANDOM}};
  regs_1201 = _RAND_1201[31:0];
  _RAND_1202 = {1{`RANDOM}};
  regs_1202 = _RAND_1202[31:0];
  _RAND_1203 = {1{`RANDOM}};
  regs_1203 = _RAND_1203[31:0];
  _RAND_1204 = {1{`RANDOM}};
  regs_1204 = _RAND_1204[31:0];
  _RAND_1205 = {1{`RANDOM}};
  regs_1205 = _RAND_1205[31:0];
  _RAND_1206 = {1{`RANDOM}};
  regs_1206 = _RAND_1206[31:0];
  _RAND_1207 = {1{`RANDOM}};
  regs_1207 = _RAND_1207[31:0];
  _RAND_1208 = {1{`RANDOM}};
  regs_1208 = _RAND_1208[31:0];
  _RAND_1209 = {1{`RANDOM}};
  regs_1209 = _RAND_1209[31:0];
  _RAND_1210 = {1{`RANDOM}};
  regs_1210 = _RAND_1210[31:0];
  _RAND_1211 = {1{`RANDOM}};
  regs_1211 = _RAND_1211[31:0];
  _RAND_1212 = {1{`RANDOM}};
  regs_1212 = _RAND_1212[31:0];
  _RAND_1213 = {1{`RANDOM}};
  regs_1213 = _RAND_1213[31:0];
  _RAND_1214 = {1{`RANDOM}};
  regs_1214 = _RAND_1214[31:0];
  _RAND_1215 = {1{`RANDOM}};
  regs_1215 = _RAND_1215[31:0];
  _RAND_1216 = {1{`RANDOM}};
  regs_1216 = _RAND_1216[31:0];
  _RAND_1217 = {1{`RANDOM}};
  regs_1217 = _RAND_1217[31:0];
  _RAND_1218 = {1{`RANDOM}};
  regs_1218 = _RAND_1218[31:0];
  _RAND_1219 = {1{`RANDOM}};
  regs_1219 = _RAND_1219[31:0];
  _RAND_1220 = {1{`RANDOM}};
  regs_1220 = _RAND_1220[31:0];
  _RAND_1221 = {1{`RANDOM}};
  regs_1221 = _RAND_1221[31:0];
  _RAND_1222 = {1{`RANDOM}};
  regs_1222 = _RAND_1222[31:0];
  _RAND_1223 = {1{`RANDOM}};
  regs_1223 = _RAND_1223[31:0];
  _RAND_1224 = {1{`RANDOM}};
  regs_1224 = _RAND_1224[31:0];
  _RAND_1225 = {1{`RANDOM}};
  regs_1225 = _RAND_1225[31:0];
  _RAND_1226 = {1{`RANDOM}};
  regs_1226 = _RAND_1226[31:0];
  _RAND_1227 = {1{`RANDOM}};
  regs_1227 = _RAND_1227[31:0];
  _RAND_1228 = {1{`RANDOM}};
  regs_1228 = _RAND_1228[31:0];
  _RAND_1229 = {1{`RANDOM}};
  regs_1229 = _RAND_1229[31:0];
  _RAND_1230 = {1{`RANDOM}};
  regs_1230 = _RAND_1230[31:0];
  _RAND_1231 = {1{`RANDOM}};
  regs_1231 = _RAND_1231[31:0];
  _RAND_1232 = {1{`RANDOM}};
  regs_1232 = _RAND_1232[31:0];
  _RAND_1233 = {1{`RANDOM}};
  regs_1233 = _RAND_1233[31:0];
  _RAND_1234 = {1{`RANDOM}};
  regs_1234 = _RAND_1234[31:0];
  _RAND_1235 = {1{`RANDOM}};
  regs_1235 = _RAND_1235[31:0];
  _RAND_1236 = {1{`RANDOM}};
  regs_1236 = _RAND_1236[31:0];
  _RAND_1237 = {1{`RANDOM}};
  regs_1237 = _RAND_1237[31:0];
  _RAND_1238 = {1{`RANDOM}};
  regs_1238 = _RAND_1238[31:0];
  _RAND_1239 = {1{`RANDOM}};
  regs_1239 = _RAND_1239[31:0];
  _RAND_1240 = {1{`RANDOM}};
  regs_1240 = _RAND_1240[31:0];
  _RAND_1241 = {1{`RANDOM}};
  regs_1241 = _RAND_1241[31:0];
  _RAND_1242 = {1{`RANDOM}};
  regs_1242 = _RAND_1242[31:0];
  _RAND_1243 = {1{`RANDOM}};
  regs_1243 = _RAND_1243[31:0];
  _RAND_1244 = {1{`RANDOM}};
  regs_1244 = _RAND_1244[31:0];
  _RAND_1245 = {1{`RANDOM}};
  regs_1245 = _RAND_1245[31:0];
  _RAND_1246 = {1{`RANDOM}};
  regs_1246 = _RAND_1246[31:0];
  _RAND_1247 = {1{`RANDOM}};
  regs_1247 = _RAND_1247[31:0];
  _RAND_1248 = {1{`RANDOM}};
  regs_1248 = _RAND_1248[31:0];
  _RAND_1249 = {1{`RANDOM}};
  regs_1249 = _RAND_1249[31:0];
  _RAND_1250 = {1{`RANDOM}};
  regs_1250 = _RAND_1250[31:0];
  _RAND_1251 = {1{`RANDOM}};
  regs_1251 = _RAND_1251[31:0];
  _RAND_1252 = {1{`RANDOM}};
  regs_1252 = _RAND_1252[31:0];
  _RAND_1253 = {1{`RANDOM}};
  regs_1253 = _RAND_1253[31:0];
  _RAND_1254 = {1{`RANDOM}};
  regs_1254 = _RAND_1254[31:0];
  _RAND_1255 = {1{`RANDOM}};
  regs_1255 = _RAND_1255[31:0];
  _RAND_1256 = {1{`RANDOM}};
  regs_1256 = _RAND_1256[31:0];
  _RAND_1257 = {1{`RANDOM}};
  regs_1257 = _RAND_1257[31:0];
  _RAND_1258 = {1{`RANDOM}};
  regs_1258 = _RAND_1258[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FP_square_root_newfpu(
  input         clock,
  input         reset,
  input         io_in_en,
  input  [31:0] io_in_a,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
`endif // RANDOMIZE_REG_INIT
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_1_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_1_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_1_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_1_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_1_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_2_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_2_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_2_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_2_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_2_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_3_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_3_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_3_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_3_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_3_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_4_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_4_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_4_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_4_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_4_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_5_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_5_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_5_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_5_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_5_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_6_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_6_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_6_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_6_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_6_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_7_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_7_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_7_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_7_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_7_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_8_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_8_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_8_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_8_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_8_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_8_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_9_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_9_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_9_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_9_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_9_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_9_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_10_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_10_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_10_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_10_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_10_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_10_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_11_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_11_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_11_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_11_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_11_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_11_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_12_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_12_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_12_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_12_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_12_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_12_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_13_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_13_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_13_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_13_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_13_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_13_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_14_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_14_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_14_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_14_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_14_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_14_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_15_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_15_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_15_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_15_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_15_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_15_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_16_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_16_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_16_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_16_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_16_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_16_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_17_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_17_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_17_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_17_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_17_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_17_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_18_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_18_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_18_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_18_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_18_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_18_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_19_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_19_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_19_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_19_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_19_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_19_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_20_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_20_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_20_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_20_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_20_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_20_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_21_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_21_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_21_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_21_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_21_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_21_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_22_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_22_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_22_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_22_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_22_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_22_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_23_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_23_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_23_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_23_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_23_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_23_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_24_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_24_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_24_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_24_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_24_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_24_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_25_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_25_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_25_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_25_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_25_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_25_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_26_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_26_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_26_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_26_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_26_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_26_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_27_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_27_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_27_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_27_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_27_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_27_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_28_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_28_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_28_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_28_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_28_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_28_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_29_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_29_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_29_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_29_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_29_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_29_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_30_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_30_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_30_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_30_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_30_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_30_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_31_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_31_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_31_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_31_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_31_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_31_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_32_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_32_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_32_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_32_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_32_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_32_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_33_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_33_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_33_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_33_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_33_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_33_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_34_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_34_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_34_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_34_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_34_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_34_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_35_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_35_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_35_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_35_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_35_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_35_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_36_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_36_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_36_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_36_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_36_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_36_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_37_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_37_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_37_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_37_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_37_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_37_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_38_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_38_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_38_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_38_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_38_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_38_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_39_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_39_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_39_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_39_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_39_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_39_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_40_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_40_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_40_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_40_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_40_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_40_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_41_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_41_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_41_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_41_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_41_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_41_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_42_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_42_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_42_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_42_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_42_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_42_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_43_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_43_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_43_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_43_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_43_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_43_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_44_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_44_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_44_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_44_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_44_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_44_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_45_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_45_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_45_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_45_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_45_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_45_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_46_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_46_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_46_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_46_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_46_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_46_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_47_clock; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_47_reset; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_multiplier_10ccs_47_io_in_en; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_47_io_in_a; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_47_io_in_b; // @[FloatingPointDesigns.scala 1985:65]
  wire [31:0] FP_multiplier_10ccs_47_io_out_s; // @[FloatingPointDesigns.scala 1985:65]
  wire  FP_subtractor_13ccs_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_1_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_1_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_1_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_1_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_1_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_2_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_2_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_2_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_2_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_2_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_3_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_3_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_3_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_3_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_3_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_3_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_4_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_4_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_4_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_4_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_4_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_4_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_5_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_5_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_5_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_5_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_5_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_5_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_6_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_6_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_6_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_6_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_6_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_6_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_7_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_7_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_7_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_7_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_7_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_7_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_8_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_8_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_8_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_8_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_8_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_8_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_9_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_9_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_9_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_9_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_9_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_9_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_10_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_10_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_10_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_10_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_10_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_10_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_11_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_11_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_11_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_11_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_11_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_11_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_12_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_12_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_12_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_12_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_12_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_12_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_13_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_13_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_13_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_13_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_13_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_13_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_14_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_14_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_14_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_14_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_14_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_14_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_15_clock; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_15_reset; // @[FloatingPointDesigns.scala 1986:50]
  wire  FP_subtractor_13ccs_15_io_in_en; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_15_io_in_a; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_15_io_in_b; // @[FloatingPointDesigns.scala 1986:50]
  wire [31:0] FP_subtractor_13ccs_15_io_out_s; // @[FloatingPointDesigns.scala 1986:50]
  wire  multiplier4_clock; // @[FloatingPointDesigns.scala 2054:29]
  wire  multiplier4_reset; // @[FloatingPointDesigns.scala 2054:29]
  wire  multiplier4_io_in_en; // @[FloatingPointDesigns.scala 2054:29]
  wire [31:0] multiplier4_io_in_a; // @[FloatingPointDesigns.scala 2054:29]
  wire [31:0] multiplier4_io_in_b; // @[FloatingPointDesigns.scala 2054:29]
  wire [31:0] multiplier4_io_out_s; // @[FloatingPointDesigns.scala 2054:29]
  wire [30:0] _number_T_1 = {{1'd0}, io_in_a[30:1]}; // @[FloatingPointDesigns.scala 1969:36]
  wire [30:0] _GEN_0 = io_in_a[30:0] > 31'h7ef477d4 ? 31'h3f7a3bea : _number_T_1; // @[FloatingPointDesigns.scala 1966:46 1967:14 1969:14]
  wire [31:0] number = {{1'd0}, _GEN_0}; // @[FloatingPointDesigns.scala 1963:22]
  wire [31:0] result = 32'h5f3759df - number; // @[FloatingPointDesigns.scala 1976:25]
  reg [31:0] x_n_0; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_1; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_2; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_4; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_5; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_6; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_8; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_9; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_10; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_12; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_13; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_14; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_16; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_17; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_18; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_20; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_21; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_22; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_24; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_25; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_26; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_28; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_29; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_30; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_32; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_33; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_34; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_36; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_37; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_38; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_40; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_41; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_42; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_44; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_45; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_46; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_48; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_49; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_50; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_52; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_53; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_54; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_56; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_57; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_58; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_60; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_61; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] x_n_62; // @[FloatingPointDesigns.scala 1978:22]
  reg [31:0] a_2_0; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_1; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_2; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_3; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_4; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_5; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_6; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_7; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_8; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_9; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_10; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_11; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_12; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_13; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_14; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_15; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_16; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_17; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_18; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_19; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_20; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_21; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_22; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_23; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_24; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_25; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_26; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_27; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_28; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_29; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_30; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_31; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_32; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_33; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_34; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_35; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_36; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_37; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_38; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_39; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_40; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_41; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_42; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_43; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_44; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_45; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_46; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_47; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_48; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_49; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_50; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_51; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_52; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_53; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_54; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_55; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_56; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_57; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_58; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_59; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_60; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_61; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_62; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] a_2_63; // @[FloatingPointDesigns.scala 1979:22]
  reg [31:0] stage1_regs_0_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_0_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_1_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_2_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_3_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_4_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_5_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_6_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_7_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_8_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_9_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_10_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_11_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_12_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_13_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_14_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_0_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_0_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_0_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_0_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_0_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_0_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_0_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_0_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_0_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_1_0; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_1_1; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_1_2; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_1_3; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_1_4; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_1_5; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_1_6; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_1_7; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage1_regs_15_1_8; // @[FloatingPointDesigns.scala 1980:30]
  reg [31:0] stage2_regs_0_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_0_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_1_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_2_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_3_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_4_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_5_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_6_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_7_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_8_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_9_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_10_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_11_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_12_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_13_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_14_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_0_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_0_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_0_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_0_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_0_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_0_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_0_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_0_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_0_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_1_0; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_1_1; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_1_2; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_1_3; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_1_4; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_1_5; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_1_6; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_1_7; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage2_regs_15_1_8; // @[FloatingPointDesigns.scala 1981:30]
  reg [31:0] stage3_regs_0_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_0_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_1_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_2_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_3_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_4_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_5_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_6_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_7_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_8_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_9_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_10_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_11_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_12_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_13_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_14_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_0_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_0_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_0_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_0_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_0_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_0_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_0_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_0_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_0_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_0_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_0_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_0_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_1_0; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_1_1; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_1_2; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_1_3; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_1_4; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_1_5; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_1_6; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_1_7; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_1_8; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_1_9; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_1_10; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage3_regs_15_1_11; // @[FloatingPointDesigns.scala 1982:30]
  reg [31:0] stage4_regs_0_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_0_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_0_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_0_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_0_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_0_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_0_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_0_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_0_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_1_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_1_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_1_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_1_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_1_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_1_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_1_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_1_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_1_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_2_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_2_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_2_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_2_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_2_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_2_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_2_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_2_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_2_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_3_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_3_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_3_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_3_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_3_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_3_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_3_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_3_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_3_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_4_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_4_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_4_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_4_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_4_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_4_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_4_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_4_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_4_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_5_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_5_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_5_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_5_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_5_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_5_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_5_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_5_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_5_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_6_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_6_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_6_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_6_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_6_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_6_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_6_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_6_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_6_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_7_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_7_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_7_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_7_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_7_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_7_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_7_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_7_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_7_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_8_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_8_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_8_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_8_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_8_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_8_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_8_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_8_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_8_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_9_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_9_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_9_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_9_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_9_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_9_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_9_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_9_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_9_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_10_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_10_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_10_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_10_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_10_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_10_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_10_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_10_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_10_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_11_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_11_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_11_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_11_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_11_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_11_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_11_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_11_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_11_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_12_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_12_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_12_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_12_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_12_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_12_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_12_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_12_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_12_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_13_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_13_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_13_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_13_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_13_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_13_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_13_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_13_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_13_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_14_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_14_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_14_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_14_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_14_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_14_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_14_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_14_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_14_1_8; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_15_1_0; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_15_1_1; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_15_1_2; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_15_1_3; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_15_1_4; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_15_1_5; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_15_1_6; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_15_1_7; // @[FloatingPointDesigns.scala 1983:30]
  reg [31:0] stage4_regs_15_1_8; // @[FloatingPointDesigns.scala 1983:30]
  wire [7:0] _a_2_0_T_3 = io_in_a[30:23] - 8'h1; // @[FloatingPointDesigns.scala 2008:75]
  wire [31:0] _a_2_0_T_6 = {io_in_a[31],_a_2_0_T_3,io_in_a[22:0]}; // @[FloatingPointDesigns.scala 2008:82]
  wire [7:0] _restore_a_T_3 = stage4_regs_15_1_8[30:23] + 8'h1; // @[FloatingPointDesigns.scala 2053:106]
  wire [8:0] _restore_a_T_4 = {stage4_regs_15_1_8[31],_restore_a_T_3}; // @[FloatingPointDesigns.scala 2053:55]
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_en(FP_multiplier_10ccs_io_in_en),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_1 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_1_clock),
    .reset(FP_multiplier_10ccs_1_reset),
    .io_in_en(FP_multiplier_10ccs_1_io_in_en),
    .io_in_a(FP_multiplier_10ccs_1_io_in_a),
    .io_in_b(FP_multiplier_10ccs_1_io_in_b),
    .io_out_s(FP_multiplier_10ccs_1_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_2 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_2_clock),
    .reset(FP_multiplier_10ccs_2_reset),
    .io_in_en(FP_multiplier_10ccs_2_io_in_en),
    .io_in_a(FP_multiplier_10ccs_2_io_in_a),
    .io_in_b(FP_multiplier_10ccs_2_io_in_b),
    .io_out_s(FP_multiplier_10ccs_2_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_3 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_3_clock),
    .reset(FP_multiplier_10ccs_3_reset),
    .io_in_en(FP_multiplier_10ccs_3_io_in_en),
    .io_in_a(FP_multiplier_10ccs_3_io_in_a),
    .io_in_b(FP_multiplier_10ccs_3_io_in_b),
    .io_out_s(FP_multiplier_10ccs_3_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_4 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_4_clock),
    .reset(FP_multiplier_10ccs_4_reset),
    .io_in_en(FP_multiplier_10ccs_4_io_in_en),
    .io_in_a(FP_multiplier_10ccs_4_io_in_a),
    .io_in_b(FP_multiplier_10ccs_4_io_in_b),
    .io_out_s(FP_multiplier_10ccs_4_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_5 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_5_clock),
    .reset(FP_multiplier_10ccs_5_reset),
    .io_in_en(FP_multiplier_10ccs_5_io_in_en),
    .io_in_a(FP_multiplier_10ccs_5_io_in_a),
    .io_in_b(FP_multiplier_10ccs_5_io_in_b),
    .io_out_s(FP_multiplier_10ccs_5_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_6 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_6_clock),
    .reset(FP_multiplier_10ccs_6_reset),
    .io_in_en(FP_multiplier_10ccs_6_io_in_en),
    .io_in_a(FP_multiplier_10ccs_6_io_in_a),
    .io_in_b(FP_multiplier_10ccs_6_io_in_b),
    .io_out_s(FP_multiplier_10ccs_6_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_7 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_7_clock),
    .reset(FP_multiplier_10ccs_7_reset),
    .io_in_en(FP_multiplier_10ccs_7_io_in_en),
    .io_in_a(FP_multiplier_10ccs_7_io_in_a),
    .io_in_b(FP_multiplier_10ccs_7_io_in_b),
    .io_out_s(FP_multiplier_10ccs_7_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_8 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_8_clock),
    .reset(FP_multiplier_10ccs_8_reset),
    .io_in_en(FP_multiplier_10ccs_8_io_in_en),
    .io_in_a(FP_multiplier_10ccs_8_io_in_a),
    .io_in_b(FP_multiplier_10ccs_8_io_in_b),
    .io_out_s(FP_multiplier_10ccs_8_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_9 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_9_clock),
    .reset(FP_multiplier_10ccs_9_reset),
    .io_in_en(FP_multiplier_10ccs_9_io_in_en),
    .io_in_a(FP_multiplier_10ccs_9_io_in_a),
    .io_in_b(FP_multiplier_10ccs_9_io_in_b),
    .io_out_s(FP_multiplier_10ccs_9_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_10 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_10_clock),
    .reset(FP_multiplier_10ccs_10_reset),
    .io_in_en(FP_multiplier_10ccs_10_io_in_en),
    .io_in_a(FP_multiplier_10ccs_10_io_in_a),
    .io_in_b(FP_multiplier_10ccs_10_io_in_b),
    .io_out_s(FP_multiplier_10ccs_10_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_11 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_11_clock),
    .reset(FP_multiplier_10ccs_11_reset),
    .io_in_en(FP_multiplier_10ccs_11_io_in_en),
    .io_in_a(FP_multiplier_10ccs_11_io_in_a),
    .io_in_b(FP_multiplier_10ccs_11_io_in_b),
    .io_out_s(FP_multiplier_10ccs_11_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_12 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_12_clock),
    .reset(FP_multiplier_10ccs_12_reset),
    .io_in_en(FP_multiplier_10ccs_12_io_in_en),
    .io_in_a(FP_multiplier_10ccs_12_io_in_a),
    .io_in_b(FP_multiplier_10ccs_12_io_in_b),
    .io_out_s(FP_multiplier_10ccs_12_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_13 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_13_clock),
    .reset(FP_multiplier_10ccs_13_reset),
    .io_in_en(FP_multiplier_10ccs_13_io_in_en),
    .io_in_a(FP_multiplier_10ccs_13_io_in_a),
    .io_in_b(FP_multiplier_10ccs_13_io_in_b),
    .io_out_s(FP_multiplier_10ccs_13_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_14 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_14_clock),
    .reset(FP_multiplier_10ccs_14_reset),
    .io_in_en(FP_multiplier_10ccs_14_io_in_en),
    .io_in_a(FP_multiplier_10ccs_14_io_in_a),
    .io_in_b(FP_multiplier_10ccs_14_io_in_b),
    .io_out_s(FP_multiplier_10ccs_14_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_15 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_15_clock),
    .reset(FP_multiplier_10ccs_15_reset),
    .io_in_en(FP_multiplier_10ccs_15_io_in_en),
    .io_in_a(FP_multiplier_10ccs_15_io_in_a),
    .io_in_b(FP_multiplier_10ccs_15_io_in_b),
    .io_out_s(FP_multiplier_10ccs_15_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_16 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_16_clock),
    .reset(FP_multiplier_10ccs_16_reset),
    .io_in_en(FP_multiplier_10ccs_16_io_in_en),
    .io_in_a(FP_multiplier_10ccs_16_io_in_a),
    .io_in_b(FP_multiplier_10ccs_16_io_in_b),
    .io_out_s(FP_multiplier_10ccs_16_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_17 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_17_clock),
    .reset(FP_multiplier_10ccs_17_reset),
    .io_in_en(FP_multiplier_10ccs_17_io_in_en),
    .io_in_a(FP_multiplier_10ccs_17_io_in_a),
    .io_in_b(FP_multiplier_10ccs_17_io_in_b),
    .io_out_s(FP_multiplier_10ccs_17_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_18 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_18_clock),
    .reset(FP_multiplier_10ccs_18_reset),
    .io_in_en(FP_multiplier_10ccs_18_io_in_en),
    .io_in_a(FP_multiplier_10ccs_18_io_in_a),
    .io_in_b(FP_multiplier_10ccs_18_io_in_b),
    .io_out_s(FP_multiplier_10ccs_18_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_19 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_19_clock),
    .reset(FP_multiplier_10ccs_19_reset),
    .io_in_en(FP_multiplier_10ccs_19_io_in_en),
    .io_in_a(FP_multiplier_10ccs_19_io_in_a),
    .io_in_b(FP_multiplier_10ccs_19_io_in_b),
    .io_out_s(FP_multiplier_10ccs_19_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_20 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_20_clock),
    .reset(FP_multiplier_10ccs_20_reset),
    .io_in_en(FP_multiplier_10ccs_20_io_in_en),
    .io_in_a(FP_multiplier_10ccs_20_io_in_a),
    .io_in_b(FP_multiplier_10ccs_20_io_in_b),
    .io_out_s(FP_multiplier_10ccs_20_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_21 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_21_clock),
    .reset(FP_multiplier_10ccs_21_reset),
    .io_in_en(FP_multiplier_10ccs_21_io_in_en),
    .io_in_a(FP_multiplier_10ccs_21_io_in_a),
    .io_in_b(FP_multiplier_10ccs_21_io_in_b),
    .io_out_s(FP_multiplier_10ccs_21_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_22 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_22_clock),
    .reset(FP_multiplier_10ccs_22_reset),
    .io_in_en(FP_multiplier_10ccs_22_io_in_en),
    .io_in_a(FP_multiplier_10ccs_22_io_in_a),
    .io_in_b(FP_multiplier_10ccs_22_io_in_b),
    .io_out_s(FP_multiplier_10ccs_22_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_23 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_23_clock),
    .reset(FP_multiplier_10ccs_23_reset),
    .io_in_en(FP_multiplier_10ccs_23_io_in_en),
    .io_in_a(FP_multiplier_10ccs_23_io_in_a),
    .io_in_b(FP_multiplier_10ccs_23_io_in_b),
    .io_out_s(FP_multiplier_10ccs_23_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_24 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_24_clock),
    .reset(FP_multiplier_10ccs_24_reset),
    .io_in_en(FP_multiplier_10ccs_24_io_in_en),
    .io_in_a(FP_multiplier_10ccs_24_io_in_a),
    .io_in_b(FP_multiplier_10ccs_24_io_in_b),
    .io_out_s(FP_multiplier_10ccs_24_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_25 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_25_clock),
    .reset(FP_multiplier_10ccs_25_reset),
    .io_in_en(FP_multiplier_10ccs_25_io_in_en),
    .io_in_a(FP_multiplier_10ccs_25_io_in_a),
    .io_in_b(FP_multiplier_10ccs_25_io_in_b),
    .io_out_s(FP_multiplier_10ccs_25_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_26 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_26_clock),
    .reset(FP_multiplier_10ccs_26_reset),
    .io_in_en(FP_multiplier_10ccs_26_io_in_en),
    .io_in_a(FP_multiplier_10ccs_26_io_in_a),
    .io_in_b(FP_multiplier_10ccs_26_io_in_b),
    .io_out_s(FP_multiplier_10ccs_26_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_27 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_27_clock),
    .reset(FP_multiplier_10ccs_27_reset),
    .io_in_en(FP_multiplier_10ccs_27_io_in_en),
    .io_in_a(FP_multiplier_10ccs_27_io_in_a),
    .io_in_b(FP_multiplier_10ccs_27_io_in_b),
    .io_out_s(FP_multiplier_10ccs_27_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_28 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_28_clock),
    .reset(FP_multiplier_10ccs_28_reset),
    .io_in_en(FP_multiplier_10ccs_28_io_in_en),
    .io_in_a(FP_multiplier_10ccs_28_io_in_a),
    .io_in_b(FP_multiplier_10ccs_28_io_in_b),
    .io_out_s(FP_multiplier_10ccs_28_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_29 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_29_clock),
    .reset(FP_multiplier_10ccs_29_reset),
    .io_in_en(FP_multiplier_10ccs_29_io_in_en),
    .io_in_a(FP_multiplier_10ccs_29_io_in_a),
    .io_in_b(FP_multiplier_10ccs_29_io_in_b),
    .io_out_s(FP_multiplier_10ccs_29_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_30 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_30_clock),
    .reset(FP_multiplier_10ccs_30_reset),
    .io_in_en(FP_multiplier_10ccs_30_io_in_en),
    .io_in_a(FP_multiplier_10ccs_30_io_in_a),
    .io_in_b(FP_multiplier_10ccs_30_io_in_b),
    .io_out_s(FP_multiplier_10ccs_30_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_31 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_31_clock),
    .reset(FP_multiplier_10ccs_31_reset),
    .io_in_en(FP_multiplier_10ccs_31_io_in_en),
    .io_in_a(FP_multiplier_10ccs_31_io_in_a),
    .io_in_b(FP_multiplier_10ccs_31_io_in_b),
    .io_out_s(FP_multiplier_10ccs_31_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_32 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_32_clock),
    .reset(FP_multiplier_10ccs_32_reset),
    .io_in_en(FP_multiplier_10ccs_32_io_in_en),
    .io_in_a(FP_multiplier_10ccs_32_io_in_a),
    .io_in_b(FP_multiplier_10ccs_32_io_in_b),
    .io_out_s(FP_multiplier_10ccs_32_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_33 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_33_clock),
    .reset(FP_multiplier_10ccs_33_reset),
    .io_in_en(FP_multiplier_10ccs_33_io_in_en),
    .io_in_a(FP_multiplier_10ccs_33_io_in_a),
    .io_in_b(FP_multiplier_10ccs_33_io_in_b),
    .io_out_s(FP_multiplier_10ccs_33_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_34 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_34_clock),
    .reset(FP_multiplier_10ccs_34_reset),
    .io_in_en(FP_multiplier_10ccs_34_io_in_en),
    .io_in_a(FP_multiplier_10ccs_34_io_in_a),
    .io_in_b(FP_multiplier_10ccs_34_io_in_b),
    .io_out_s(FP_multiplier_10ccs_34_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_35 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_35_clock),
    .reset(FP_multiplier_10ccs_35_reset),
    .io_in_en(FP_multiplier_10ccs_35_io_in_en),
    .io_in_a(FP_multiplier_10ccs_35_io_in_a),
    .io_in_b(FP_multiplier_10ccs_35_io_in_b),
    .io_out_s(FP_multiplier_10ccs_35_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_36 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_36_clock),
    .reset(FP_multiplier_10ccs_36_reset),
    .io_in_en(FP_multiplier_10ccs_36_io_in_en),
    .io_in_a(FP_multiplier_10ccs_36_io_in_a),
    .io_in_b(FP_multiplier_10ccs_36_io_in_b),
    .io_out_s(FP_multiplier_10ccs_36_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_37 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_37_clock),
    .reset(FP_multiplier_10ccs_37_reset),
    .io_in_en(FP_multiplier_10ccs_37_io_in_en),
    .io_in_a(FP_multiplier_10ccs_37_io_in_a),
    .io_in_b(FP_multiplier_10ccs_37_io_in_b),
    .io_out_s(FP_multiplier_10ccs_37_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_38 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_38_clock),
    .reset(FP_multiplier_10ccs_38_reset),
    .io_in_en(FP_multiplier_10ccs_38_io_in_en),
    .io_in_a(FP_multiplier_10ccs_38_io_in_a),
    .io_in_b(FP_multiplier_10ccs_38_io_in_b),
    .io_out_s(FP_multiplier_10ccs_38_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_39 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_39_clock),
    .reset(FP_multiplier_10ccs_39_reset),
    .io_in_en(FP_multiplier_10ccs_39_io_in_en),
    .io_in_a(FP_multiplier_10ccs_39_io_in_a),
    .io_in_b(FP_multiplier_10ccs_39_io_in_b),
    .io_out_s(FP_multiplier_10ccs_39_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_40 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_40_clock),
    .reset(FP_multiplier_10ccs_40_reset),
    .io_in_en(FP_multiplier_10ccs_40_io_in_en),
    .io_in_a(FP_multiplier_10ccs_40_io_in_a),
    .io_in_b(FP_multiplier_10ccs_40_io_in_b),
    .io_out_s(FP_multiplier_10ccs_40_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_41 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_41_clock),
    .reset(FP_multiplier_10ccs_41_reset),
    .io_in_en(FP_multiplier_10ccs_41_io_in_en),
    .io_in_a(FP_multiplier_10ccs_41_io_in_a),
    .io_in_b(FP_multiplier_10ccs_41_io_in_b),
    .io_out_s(FP_multiplier_10ccs_41_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_42 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_42_clock),
    .reset(FP_multiplier_10ccs_42_reset),
    .io_in_en(FP_multiplier_10ccs_42_io_in_en),
    .io_in_a(FP_multiplier_10ccs_42_io_in_a),
    .io_in_b(FP_multiplier_10ccs_42_io_in_b),
    .io_out_s(FP_multiplier_10ccs_42_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_43 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_43_clock),
    .reset(FP_multiplier_10ccs_43_reset),
    .io_in_en(FP_multiplier_10ccs_43_io_in_en),
    .io_in_a(FP_multiplier_10ccs_43_io_in_a),
    .io_in_b(FP_multiplier_10ccs_43_io_in_b),
    .io_out_s(FP_multiplier_10ccs_43_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_44 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_44_clock),
    .reset(FP_multiplier_10ccs_44_reset),
    .io_in_en(FP_multiplier_10ccs_44_io_in_en),
    .io_in_a(FP_multiplier_10ccs_44_io_in_a),
    .io_in_b(FP_multiplier_10ccs_44_io_in_b),
    .io_out_s(FP_multiplier_10ccs_44_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_45 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_45_clock),
    .reset(FP_multiplier_10ccs_45_reset),
    .io_in_en(FP_multiplier_10ccs_45_io_in_en),
    .io_in_a(FP_multiplier_10ccs_45_io_in_a),
    .io_in_b(FP_multiplier_10ccs_45_io_in_b),
    .io_out_s(FP_multiplier_10ccs_45_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_46 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_46_clock),
    .reset(FP_multiplier_10ccs_46_reset),
    .io_in_en(FP_multiplier_10ccs_46_io_in_en),
    .io_in_a(FP_multiplier_10ccs_46_io_in_a),
    .io_in_b(FP_multiplier_10ccs_46_io_in_b),
    .io_out_s(FP_multiplier_10ccs_46_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_47 ( // @[FloatingPointDesigns.scala 1985:65]
    .clock(FP_multiplier_10ccs_47_clock),
    .reset(FP_multiplier_10ccs_47_reset),
    .io_in_en(FP_multiplier_10ccs_47_io_in_en),
    .io_in_a(FP_multiplier_10ccs_47_io_in_a),
    .io_in_b(FP_multiplier_10ccs_47_io_in_b),
    .io_out_s(FP_multiplier_10ccs_47_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_clock),
    .reset(FP_subtractor_13ccs_reset),
    .io_in_en(FP_subtractor_13ccs_io_in_en),
    .io_in_a(FP_subtractor_13ccs_io_in_a),
    .io_in_b(FP_subtractor_13ccs_io_in_b),
    .io_out_s(FP_subtractor_13ccs_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_1 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_1_clock),
    .reset(FP_subtractor_13ccs_1_reset),
    .io_in_en(FP_subtractor_13ccs_1_io_in_en),
    .io_in_a(FP_subtractor_13ccs_1_io_in_a),
    .io_in_b(FP_subtractor_13ccs_1_io_in_b),
    .io_out_s(FP_subtractor_13ccs_1_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_2 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_2_clock),
    .reset(FP_subtractor_13ccs_2_reset),
    .io_in_en(FP_subtractor_13ccs_2_io_in_en),
    .io_in_a(FP_subtractor_13ccs_2_io_in_a),
    .io_in_b(FP_subtractor_13ccs_2_io_in_b),
    .io_out_s(FP_subtractor_13ccs_2_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_3 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_3_clock),
    .reset(FP_subtractor_13ccs_3_reset),
    .io_in_en(FP_subtractor_13ccs_3_io_in_en),
    .io_in_a(FP_subtractor_13ccs_3_io_in_a),
    .io_in_b(FP_subtractor_13ccs_3_io_in_b),
    .io_out_s(FP_subtractor_13ccs_3_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_4 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_4_clock),
    .reset(FP_subtractor_13ccs_4_reset),
    .io_in_en(FP_subtractor_13ccs_4_io_in_en),
    .io_in_a(FP_subtractor_13ccs_4_io_in_a),
    .io_in_b(FP_subtractor_13ccs_4_io_in_b),
    .io_out_s(FP_subtractor_13ccs_4_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_5 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_5_clock),
    .reset(FP_subtractor_13ccs_5_reset),
    .io_in_en(FP_subtractor_13ccs_5_io_in_en),
    .io_in_a(FP_subtractor_13ccs_5_io_in_a),
    .io_in_b(FP_subtractor_13ccs_5_io_in_b),
    .io_out_s(FP_subtractor_13ccs_5_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_6 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_6_clock),
    .reset(FP_subtractor_13ccs_6_reset),
    .io_in_en(FP_subtractor_13ccs_6_io_in_en),
    .io_in_a(FP_subtractor_13ccs_6_io_in_a),
    .io_in_b(FP_subtractor_13ccs_6_io_in_b),
    .io_out_s(FP_subtractor_13ccs_6_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_7 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_7_clock),
    .reset(FP_subtractor_13ccs_7_reset),
    .io_in_en(FP_subtractor_13ccs_7_io_in_en),
    .io_in_a(FP_subtractor_13ccs_7_io_in_a),
    .io_in_b(FP_subtractor_13ccs_7_io_in_b),
    .io_out_s(FP_subtractor_13ccs_7_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_8 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_8_clock),
    .reset(FP_subtractor_13ccs_8_reset),
    .io_in_en(FP_subtractor_13ccs_8_io_in_en),
    .io_in_a(FP_subtractor_13ccs_8_io_in_a),
    .io_in_b(FP_subtractor_13ccs_8_io_in_b),
    .io_out_s(FP_subtractor_13ccs_8_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_9 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_9_clock),
    .reset(FP_subtractor_13ccs_9_reset),
    .io_in_en(FP_subtractor_13ccs_9_io_in_en),
    .io_in_a(FP_subtractor_13ccs_9_io_in_a),
    .io_in_b(FP_subtractor_13ccs_9_io_in_b),
    .io_out_s(FP_subtractor_13ccs_9_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_10 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_10_clock),
    .reset(FP_subtractor_13ccs_10_reset),
    .io_in_en(FP_subtractor_13ccs_10_io_in_en),
    .io_in_a(FP_subtractor_13ccs_10_io_in_a),
    .io_in_b(FP_subtractor_13ccs_10_io_in_b),
    .io_out_s(FP_subtractor_13ccs_10_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_11 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_11_clock),
    .reset(FP_subtractor_13ccs_11_reset),
    .io_in_en(FP_subtractor_13ccs_11_io_in_en),
    .io_in_a(FP_subtractor_13ccs_11_io_in_a),
    .io_in_b(FP_subtractor_13ccs_11_io_in_b),
    .io_out_s(FP_subtractor_13ccs_11_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_12 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_12_clock),
    .reset(FP_subtractor_13ccs_12_reset),
    .io_in_en(FP_subtractor_13ccs_12_io_in_en),
    .io_in_a(FP_subtractor_13ccs_12_io_in_a),
    .io_in_b(FP_subtractor_13ccs_12_io_in_b),
    .io_out_s(FP_subtractor_13ccs_12_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_13 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_13_clock),
    .reset(FP_subtractor_13ccs_13_reset),
    .io_in_en(FP_subtractor_13ccs_13_io_in_en),
    .io_in_a(FP_subtractor_13ccs_13_io_in_a),
    .io_in_b(FP_subtractor_13ccs_13_io_in_b),
    .io_out_s(FP_subtractor_13ccs_13_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_14 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_14_clock),
    .reset(FP_subtractor_13ccs_14_reset),
    .io_in_en(FP_subtractor_13ccs_14_io_in_en),
    .io_in_a(FP_subtractor_13ccs_14_io_in_a),
    .io_in_b(FP_subtractor_13ccs_14_io_in_b),
    .io_out_s(FP_subtractor_13ccs_14_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_15 ( // @[FloatingPointDesigns.scala 1986:50]
    .clock(FP_subtractor_13ccs_15_clock),
    .reset(FP_subtractor_13ccs_15_reset),
    .io_in_en(FP_subtractor_13ccs_15_io_in_en),
    .io_in_a(FP_subtractor_13ccs_15_io_in_a),
    .io_in_b(FP_subtractor_13ccs_15_io_in_b),
    .io_out_s(FP_subtractor_13ccs_15_io_out_s)
  );
  FP_multiplier_10ccs multiplier4 ( // @[FloatingPointDesigns.scala 2054:29]
    .clock(multiplier4_clock),
    .reset(multiplier4_reset),
    .io_in_en(multiplier4_io_in_en),
    .io_in_a(multiplier4_io_in_a),
    .io_in_b(multiplier4_io_in_b),
    .io_out_s(multiplier4_io_out_s)
  );
  assign io_out_s = {{1'd0}, multiplier4_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2058:14]
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_io_in_a = {1'h0,result[30:0]}; // @[FloatingPointDesigns.scala 2012:48]
  assign FP_multiplier_10ccs_io_in_b = {1'h0,result[30:0]}; // @[FloatingPointDesigns.scala 2013:48]
  assign FP_multiplier_10ccs_1_clock = clock;
  assign FP_multiplier_10ccs_1_reset = reset;
  assign FP_multiplier_10ccs_1_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_1_io_in_a = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_1_io_in_b = {1'h0,stage1_regs_0_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_2_clock = clock;
  assign FP_multiplier_10ccs_2_reset = reset;
  assign FP_multiplier_10ccs_2_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_2_io_in_a = {1'h0,stage3_regs_0_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_2_io_in_b = FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_3_clock = clock;
  assign FP_multiplier_10ccs_3_reset = reset;
  assign FP_multiplier_10ccs_3_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_3_io_in_a = {1'h0,FP_multiplier_10ccs_2_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_3_io_in_b = {1'h0,FP_multiplier_10ccs_2_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_4_clock = clock;
  assign FP_multiplier_10ccs_4_reset = reset;
  assign FP_multiplier_10ccs_4_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_4_io_in_a = FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_4_io_in_b = {1'h0,stage1_regs_1_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_5_clock = clock;
  assign FP_multiplier_10ccs_5_reset = reset;
  assign FP_multiplier_10ccs_5_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_5_io_in_a = {1'h0,stage3_regs_1_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_5_io_in_b = FP_subtractor_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_6_clock = clock;
  assign FP_multiplier_10ccs_6_reset = reset;
  assign FP_multiplier_10ccs_6_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_6_io_in_a = {1'h0,FP_multiplier_10ccs_5_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_6_io_in_b = {1'h0,FP_multiplier_10ccs_5_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_7_clock = clock;
  assign FP_multiplier_10ccs_7_reset = reset;
  assign FP_multiplier_10ccs_7_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_7_io_in_a = FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_7_io_in_b = {1'h0,stage1_regs_2_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_8_clock = clock;
  assign FP_multiplier_10ccs_8_reset = reset;
  assign FP_multiplier_10ccs_8_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_8_io_in_a = {1'h0,stage3_regs_2_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_8_io_in_b = FP_subtractor_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_9_clock = clock;
  assign FP_multiplier_10ccs_9_reset = reset;
  assign FP_multiplier_10ccs_9_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_9_io_in_a = {1'h0,FP_multiplier_10ccs_8_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_9_io_in_b = {1'h0,FP_multiplier_10ccs_8_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_10_clock = clock;
  assign FP_multiplier_10ccs_10_reset = reset;
  assign FP_multiplier_10ccs_10_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_10_io_in_a = FP_multiplier_10ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_10_io_in_b = {1'h0,stage1_regs_3_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_11_clock = clock;
  assign FP_multiplier_10ccs_11_reset = reset;
  assign FP_multiplier_10ccs_11_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_11_io_in_a = {1'h0,stage3_regs_3_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_11_io_in_b = FP_subtractor_13ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_12_clock = clock;
  assign FP_multiplier_10ccs_12_reset = reset;
  assign FP_multiplier_10ccs_12_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_12_io_in_a = {1'h0,FP_multiplier_10ccs_11_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_12_io_in_b = {1'h0,FP_multiplier_10ccs_11_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_13_clock = clock;
  assign FP_multiplier_10ccs_13_reset = reset;
  assign FP_multiplier_10ccs_13_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_13_io_in_a = FP_multiplier_10ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_13_io_in_b = {1'h0,stage1_regs_4_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_14_clock = clock;
  assign FP_multiplier_10ccs_14_reset = reset;
  assign FP_multiplier_10ccs_14_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_14_io_in_a = {1'h0,stage3_regs_4_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_14_io_in_b = FP_subtractor_13ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_15_clock = clock;
  assign FP_multiplier_10ccs_15_reset = reset;
  assign FP_multiplier_10ccs_15_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_15_io_in_a = {1'h0,FP_multiplier_10ccs_14_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_15_io_in_b = {1'h0,FP_multiplier_10ccs_14_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_16_clock = clock;
  assign FP_multiplier_10ccs_16_reset = reset;
  assign FP_multiplier_10ccs_16_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_16_io_in_a = FP_multiplier_10ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_16_io_in_b = {1'h0,stage1_regs_5_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_17_clock = clock;
  assign FP_multiplier_10ccs_17_reset = reset;
  assign FP_multiplier_10ccs_17_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_17_io_in_a = {1'h0,stage3_regs_5_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_17_io_in_b = FP_subtractor_13ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_18_clock = clock;
  assign FP_multiplier_10ccs_18_reset = reset;
  assign FP_multiplier_10ccs_18_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_18_io_in_a = {1'h0,FP_multiplier_10ccs_17_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_18_io_in_b = {1'h0,FP_multiplier_10ccs_17_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_19_clock = clock;
  assign FP_multiplier_10ccs_19_reset = reset;
  assign FP_multiplier_10ccs_19_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_19_io_in_a = FP_multiplier_10ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_19_io_in_b = {1'h0,stage1_regs_6_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_20_clock = clock;
  assign FP_multiplier_10ccs_20_reset = reset;
  assign FP_multiplier_10ccs_20_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_20_io_in_a = {1'h0,stage3_regs_6_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_20_io_in_b = FP_subtractor_13ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_21_clock = clock;
  assign FP_multiplier_10ccs_21_reset = reset;
  assign FP_multiplier_10ccs_21_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_21_io_in_a = {1'h0,FP_multiplier_10ccs_20_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_21_io_in_b = {1'h0,FP_multiplier_10ccs_20_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_22_clock = clock;
  assign FP_multiplier_10ccs_22_reset = reset;
  assign FP_multiplier_10ccs_22_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_22_io_in_a = FP_multiplier_10ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_22_io_in_b = {1'h0,stage1_regs_7_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_23_clock = clock;
  assign FP_multiplier_10ccs_23_reset = reset;
  assign FP_multiplier_10ccs_23_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_23_io_in_a = {1'h0,stage3_regs_7_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_23_io_in_b = FP_subtractor_13ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_24_clock = clock;
  assign FP_multiplier_10ccs_24_reset = reset;
  assign FP_multiplier_10ccs_24_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_24_io_in_a = {1'h0,FP_multiplier_10ccs_23_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_24_io_in_b = {1'h0,FP_multiplier_10ccs_23_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_25_clock = clock;
  assign FP_multiplier_10ccs_25_reset = reset;
  assign FP_multiplier_10ccs_25_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_25_io_in_a = FP_multiplier_10ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_25_io_in_b = {1'h0,stage1_regs_8_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_26_clock = clock;
  assign FP_multiplier_10ccs_26_reset = reset;
  assign FP_multiplier_10ccs_26_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_26_io_in_a = {1'h0,stage3_regs_8_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_26_io_in_b = FP_subtractor_13ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_27_clock = clock;
  assign FP_multiplier_10ccs_27_reset = reset;
  assign FP_multiplier_10ccs_27_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_27_io_in_a = {1'h0,FP_multiplier_10ccs_26_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_27_io_in_b = {1'h0,FP_multiplier_10ccs_26_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_28_clock = clock;
  assign FP_multiplier_10ccs_28_reset = reset;
  assign FP_multiplier_10ccs_28_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_28_io_in_a = FP_multiplier_10ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_28_io_in_b = {1'h0,stage1_regs_9_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_29_clock = clock;
  assign FP_multiplier_10ccs_29_reset = reset;
  assign FP_multiplier_10ccs_29_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_29_io_in_a = {1'h0,stage3_regs_9_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_29_io_in_b = FP_subtractor_13ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_30_clock = clock;
  assign FP_multiplier_10ccs_30_reset = reset;
  assign FP_multiplier_10ccs_30_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_30_io_in_a = {1'h0,FP_multiplier_10ccs_29_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_30_io_in_b = {1'h0,FP_multiplier_10ccs_29_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_31_clock = clock;
  assign FP_multiplier_10ccs_31_reset = reset;
  assign FP_multiplier_10ccs_31_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_31_io_in_a = FP_multiplier_10ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_31_io_in_b = {1'h0,stage1_regs_10_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_32_clock = clock;
  assign FP_multiplier_10ccs_32_reset = reset;
  assign FP_multiplier_10ccs_32_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_32_io_in_a = {1'h0,stage3_regs_10_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_32_io_in_b = FP_subtractor_13ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_33_clock = clock;
  assign FP_multiplier_10ccs_33_reset = reset;
  assign FP_multiplier_10ccs_33_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_33_io_in_a = {1'h0,FP_multiplier_10ccs_32_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_33_io_in_b = {1'h0,FP_multiplier_10ccs_32_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_34_clock = clock;
  assign FP_multiplier_10ccs_34_reset = reset;
  assign FP_multiplier_10ccs_34_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_34_io_in_a = FP_multiplier_10ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_34_io_in_b = {1'h0,stage1_regs_11_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_35_clock = clock;
  assign FP_multiplier_10ccs_35_reset = reset;
  assign FP_multiplier_10ccs_35_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_35_io_in_a = {1'h0,stage3_regs_11_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_35_io_in_b = FP_subtractor_13ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_36_clock = clock;
  assign FP_multiplier_10ccs_36_reset = reset;
  assign FP_multiplier_10ccs_36_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_36_io_in_a = {1'h0,FP_multiplier_10ccs_35_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_36_io_in_b = {1'h0,FP_multiplier_10ccs_35_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_37_clock = clock;
  assign FP_multiplier_10ccs_37_reset = reset;
  assign FP_multiplier_10ccs_37_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_37_io_in_a = FP_multiplier_10ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_37_io_in_b = {1'h0,stage1_regs_12_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_38_clock = clock;
  assign FP_multiplier_10ccs_38_reset = reset;
  assign FP_multiplier_10ccs_38_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_38_io_in_a = {1'h0,stage3_regs_12_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_38_io_in_b = FP_subtractor_13ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_39_clock = clock;
  assign FP_multiplier_10ccs_39_reset = reset;
  assign FP_multiplier_10ccs_39_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_39_io_in_a = {1'h0,FP_multiplier_10ccs_38_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_39_io_in_b = {1'h0,FP_multiplier_10ccs_38_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_40_clock = clock;
  assign FP_multiplier_10ccs_40_reset = reset;
  assign FP_multiplier_10ccs_40_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_40_io_in_a = FP_multiplier_10ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_40_io_in_b = {1'h0,stage1_regs_13_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_41_clock = clock;
  assign FP_multiplier_10ccs_41_reset = reset;
  assign FP_multiplier_10ccs_41_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_41_io_in_a = {1'h0,stage3_regs_13_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_41_io_in_b = FP_subtractor_13ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_42_clock = clock;
  assign FP_multiplier_10ccs_42_reset = reset;
  assign FP_multiplier_10ccs_42_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_42_io_in_a = {1'h0,FP_multiplier_10ccs_41_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_42_io_in_b = {1'h0,FP_multiplier_10ccs_41_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_43_clock = clock;
  assign FP_multiplier_10ccs_43_reset = reset;
  assign FP_multiplier_10ccs_43_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_43_io_in_a = FP_multiplier_10ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_43_io_in_b = {1'h0,stage1_regs_14_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_44_clock = clock;
  assign FP_multiplier_10ccs_44_reset = reset;
  assign FP_multiplier_10ccs_44_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_44_io_in_a = {1'h0,stage3_regs_14_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_44_io_in_b = FP_subtractor_13ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_multiplier_10ccs_45_clock = clock;
  assign FP_multiplier_10ccs_45_reset = reset;
  assign FP_multiplier_10ccs_45_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_45_io_in_a = {1'h0,FP_multiplier_10ccs_44_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2021:48]
  assign FP_multiplier_10ccs_45_io_in_b = {1'h0,FP_multiplier_10ccs_44_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2022:48]
  assign FP_multiplier_10ccs_46_clock = clock;
  assign FP_multiplier_10ccs_46_reset = reset;
  assign FP_multiplier_10ccs_46_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_46_io_in_a = FP_multiplier_10ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2025:34]
  assign FP_multiplier_10ccs_46_io_in_b = {1'h0,stage1_regs_15_1_8[30:0]}; // @[FloatingPointDesigns.scala 2026:46]
  assign FP_multiplier_10ccs_47_clock = clock;
  assign FP_multiplier_10ccs_47_reset = reset;
  assign FP_multiplier_10ccs_47_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1987:41]
  assign FP_multiplier_10ccs_47_io_in_a = {1'h0,stage3_regs_15_0_11[30:0]}; // @[FloatingPointDesigns.scala 2043:46]
  assign FP_multiplier_10ccs_47_io_in_b = FP_subtractor_13ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2044:34]
  assign FP_subtractor_13ccs_clock = clock;
  assign FP_subtractor_13ccs_reset = reset;
  assign FP_subtractor_13ccs_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_io_in_b = FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_1_clock = clock;
  assign FP_subtractor_13ccs_1_reset = reset;
  assign FP_subtractor_13ccs_1_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_1_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_1_io_in_b = FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_2_clock = clock;
  assign FP_subtractor_13ccs_2_reset = reset;
  assign FP_subtractor_13ccs_2_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_2_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_2_io_in_b = FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_3_clock = clock;
  assign FP_subtractor_13ccs_3_reset = reset;
  assign FP_subtractor_13ccs_3_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_3_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_3_io_in_b = FP_multiplier_10ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_4_clock = clock;
  assign FP_subtractor_13ccs_4_reset = reset;
  assign FP_subtractor_13ccs_4_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_4_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_4_io_in_b = FP_multiplier_10ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_5_clock = clock;
  assign FP_subtractor_13ccs_5_reset = reset;
  assign FP_subtractor_13ccs_5_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_5_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_5_io_in_b = FP_multiplier_10ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_6_clock = clock;
  assign FP_subtractor_13ccs_6_reset = reset;
  assign FP_subtractor_13ccs_6_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_6_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_6_io_in_b = FP_multiplier_10ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_7_clock = clock;
  assign FP_subtractor_13ccs_7_reset = reset;
  assign FP_subtractor_13ccs_7_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_7_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_7_io_in_b = FP_multiplier_10ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_8_clock = clock;
  assign FP_subtractor_13ccs_8_reset = reset;
  assign FP_subtractor_13ccs_8_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_8_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_8_io_in_b = FP_multiplier_10ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_9_clock = clock;
  assign FP_subtractor_13ccs_9_reset = reset;
  assign FP_subtractor_13ccs_9_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_9_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_9_io_in_b = FP_multiplier_10ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_10_clock = clock;
  assign FP_subtractor_13ccs_10_reset = reset;
  assign FP_subtractor_13ccs_10_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_10_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_10_io_in_b = FP_multiplier_10ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_11_clock = clock;
  assign FP_subtractor_13ccs_11_reset = reset;
  assign FP_subtractor_13ccs_11_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_11_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_11_io_in_b = FP_multiplier_10ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_12_clock = clock;
  assign FP_subtractor_13ccs_12_reset = reset;
  assign FP_subtractor_13ccs_12_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_12_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_12_io_in_b = FP_multiplier_10ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_13_clock = clock;
  assign FP_subtractor_13ccs_13_reset = reset;
  assign FP_subtractor_13ccs_13_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_13_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_13_io_in_b = FP_multiplier_10ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_14_clock = clock;
  assign FP_subtractor_13ccs_14_reset = reset;
  assign FP_subtractor_13ccs_14_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_14_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_14_io_in_b = FP_multiplier_10ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign FP_subtractor_13ccs_15_clock = clock;
  assign FP_subtractor_13ccs_15_reset = reset;
  assign FP_subtractor_13ccs_15_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 1988:32]
  assign FP_subtractor_13ccs_15_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1964:26 1965:16]
  assign FP_subtractor_13ccs_15_io_in_b = FP_multiplier_10ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2035:31]
  assign multiplier4_clock = clock;
  assign multiplier4_reset = reset;
  assign multiplier4_io_in_en = io_in_en; // @[FloatingPointDesigns.scala 2055:26]
  assign multiplier4_io_in_a = {1'h0,FP_multiplier_10ccs_47_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2056:37]
  assign multiplier4_io_in_b = {_restore_a_T_4,stage4_regs_15_1_8[22:0]}; // @[FloatingPointDesigns.scala 2053:113]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_0 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2006:28]
      x_n_0 <= result; // @[FloatingPointDesigns.scala 2007:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_1 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_1 <= stage1_regs_0_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_2 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_2 <= stage2_regs_0_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_4 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_4 <= FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_5 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_5 <= stage1_regs_1_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_6 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_6 <= stage2_regs_1_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_8 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_8 <= FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_9 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_9 <= stage1_regs_2_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_10 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_10 <= stage2_regs_2_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_12 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_12 <= FP_multiplier_10ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_13 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_13 <= stage1_regs_3_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_14 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_14 <= stage2_regs_3_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_16 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_16 <= FP_multiplier_10ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_17 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_17 <= stage1_regs_4_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_18 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_18 <= stage2_regs_4_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_20 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_20 <= FP_multiplier_10ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_21 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_21 <= stage1_regs_5_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_22 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_22 <= stage2_regs_5_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_24 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_24 <= FP_multiplier_10ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_25 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_25 <= stage1_regs_6_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_26 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_26 <= stage2_regs_6_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_28 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_28 <= FP_multiplier_10ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_29 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_29 <= stage1_regs_7_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_30 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_30 <= stage2_regs_7_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_32 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_32 <= FP_multiplier_10ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_33 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_33 <= stage1_regs_8_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_34 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_34 <= stage2_regs_8_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_36 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_36 <= FP_multiplier_10ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_37 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_37 <= stage1_regs_9_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_38 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_38 <= stage2_regs_9_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_40 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_40 <= FP_multiplier_10ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_41 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_41 <= stage1_regs_10_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_42 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_42 <= stage2_regs_10_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_44 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_44 <= FP_multiplier_10ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_45 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_45 <= stage1_regs_11_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_46 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_46 <= stage2_regs_11_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_48 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_48 <= FP_multiplier_10ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_49 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_49 <= stage1_regs_12_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_50 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_50 <= stage2_regs_12_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_52 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_52 <= FP_multiplier_10ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_53 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_53 <= stage1_regs_13_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_54 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_54 <= stage2_regs_13_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_56 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_56 <= FP_multiplier_10ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_57 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_57 <= stage1_regs_14_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_58 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_58 <= stage2_regs_14_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_60 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      x_n_60 <= FP_multiplier_10ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2016:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_61 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      x_n_61 <= stage1_regs_15_0_8; // @[FloatingPointDesigns.scala 2029:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1978:22]
      x_n_62 <= 32'h0; // @[FloatingPointDesigns.scala 1978:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      x_n_62 <= stage2_regs_15_0_8; // @[FloatingPointDesigns.scala 2038:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_0 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2006:28]
      a_2_0 <= _a_2_0_T_6; // @[FloatingPointDesigns.scala 2008:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_1 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_1 <= stage1_regs_0_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_2 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_2 <= stage2_regs_0_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_3 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_3 <= stage3_regs_0_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_4 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_4 <= stage4_regs_0_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_5 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_5 <= stage1_regs_1_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_6 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_6 <= stage2_regs_1_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_7 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_7 <= stage3_regs_1_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_8 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_8 <= stage4_regs_1_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_9 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_9 <= stage1_regs_2_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_10 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_10 <= stage2_regs_2_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_11 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_11 <= stage3_regs_2_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_12 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_12 <= stage4_regs_2_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_13 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_13 <= stage1_regs_3_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_14 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_14 <= stage2_regs_3_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_15 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_15 <= stage3_regs_3_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_16 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_16 <= stage4_regs_3_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_17 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_17 <= stage1_regs_4_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_18 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_18 <= stage2_regs_4_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_19 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_19 <= stage3_regs_4_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_20 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_20 <= stage4_regs_4_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_21 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_21 <= stage1_regs_5_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_22 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_22 <= stage2_regs_5_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_23 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_23 <= stage3_regs_5_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_24 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_24 <= stage4_regs_5_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_25 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_25 <= stage1_regs_6_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_26 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_26 <= stage2_regs_6_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_27 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_27 <= stage3_regs_6_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_28 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_28 <= stage4_regs_6_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_29 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_29 <= stage1_regs_7_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_30 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_30 <= stage2_regs_7_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_31 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_31 <= stage3_regs_7_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_32 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_32 <= stage4_regs_7_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_33 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_33 <= stage1_regs_8_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_34 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_34 <= stage2_regs_8_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_35 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_35 <= stage3_regs_8_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_36 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_36 <= stage4_regs_8_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_37 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_37 <= stage1_regs_9_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_38 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_38 <= stage2_regs_9_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_39 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_39 <= stage3_regs_9_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_40 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_40 <= stage4_regs_9_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_41 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_41 <= stage1_regs_10_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_42 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_42 <= stage2_regs_10_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_43 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_43 <= stage3_regs_10_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_44 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_44 <= stage4_regs_10_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_45 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_45 <= stage1_regs_11_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_46 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_46 <= stage2_regs_11_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_47 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_47 <= stage3_regs_11_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_48 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_48 <= stage4_regs_11_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_49 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_49 <= stage1_regs_12_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_50 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_50 <= stage2_regs_12_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_51 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_51 <= stage3_regs_12_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_52 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_52 <= stage4_regs_12_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_53 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_53 <= stage1_regs_13_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_54 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_54 <= stage2_regs_13_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_55 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_55 <= stage3_regs_13_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_56 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_56 <= stage4_regs_13_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_57 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_57 <= stage1_regs_14_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_58 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_58 <= stage2_regs_14_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_59 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_59 <= stage3_regs_14_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_60 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      a_2_60 <= stage4_regs_14_1_8; // @[FloatingPointDesigns.scala 2017:26]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_61 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      a_2_61 <= stage1_regs_15_1_8; // @[FloatingPointDesigns.scala 2028:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_62 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      a_2_62 <= stage2_regs_15_1_8; // @[FloatingPointDesigns.scala 2037:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1979:22]
      a_2_63 <= 32'h0; // @[FloatingPointDesigns.scala 1979:22]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      a_2_63 <= stage3_regs_15_1_11; // @[FloatingPointDesigns.scala 2046:28]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2006:28]
      stage1_regs_0_0_0 <= x_n_0; // @[FloatingPointDesigns.scala 2009:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_0_1 <= stage1_regs_0_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_0_2 <= stage1_regs_0_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_0_3 <= stage1_regs_0_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_0_4 <= stage1_regs_0_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_0_5 <= stage1_regs_0_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_0_6 <= stage1_regs_0_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_0_7 <= stage1_regs_0_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_0_8 <= stage1_regs_0_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2006:28]
      stage1_regs_0_1_0 <= a_2_0; // @[FloatingPointDesigns.scala 2010:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_1_1 <= stage1_regs_0_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_1_2 <= stage1_regs_0_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_1_3 <= stage1_regs_0_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_1_4 <= stage1_regs_0_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_1_5 <= stage1_regs_0_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_1_6 <= stage1_regs_0_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_1_7 <= stage1_regs_0_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_0_1_8 <= stage1_regs_0_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_1_0_0 <= x_n_4; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_0_1 <= stage1_regs_1_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_0_2 <= stage1_regs_1_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_0_3 <= stage1_regs_1_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_0_4 <= stage1_regs_1_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_0_5 <= stage1_regs_1_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_0_6 <= stage1_regs_1_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_0_7 <= stage1_regs_1_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_0_8 <= stage1_regs_1_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_1_1_0 <= a_2_4; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_1_1 <= stage1_regs_1_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_1_2 <= stage1_regs_1_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_1_3 <= stage1_regs_1_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_1_4 <= stage1_regs_1_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_1_5 <= stage1_regs_1_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_1_6 <= stage1_regs_1_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_1_7 <= stage1_regs_1_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_1_1_8 <= stage1_regs_1_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_2_0_0 <= x_n_8; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_0_1 <= stage1_regs_2_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_0_2 <= stage1_regs_2_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_0_3 <= stage1_regs_2_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_0_4 <= stage1_regs_2_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_0_5 <= stage1_regs_2_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_0_6 <= stage1_regs_2_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_0_7 <= stage1_regs_2_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_0_8 <= stage1_regs_2_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_2_1_0 <= a_2_8; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_1_1 <= stage1_regs_2_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_1_2 <= stage1_regs_2_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_1_3 <= stage1_regs_2_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_1_4 <= stage1_regs_2_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_1_5 <= stage1_regs_2_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_1_6 <= stage1_regs_2_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_1_7 <= stage1_regs_2_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_2_1_8 <= stage1_regs_2_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_3_0_0 <= x_n_12; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_0_1 <= stage1_regs_3_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_0_2 <= stage1_regs_3_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_0_3 <= stage1_regs_3_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_0_4 <= stage1_regs_3_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_0_5 <= stage1_regs_3_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_0_6 <= stage1_regs_3_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_0_7 <= stage1_regs_3_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_0_8 <= stage1_regs_3_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_3_1_0 <= a_2_12; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_1_1 <= stage1_regs_3_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_1_2 <= stage1_regs_3_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_1_3 <= stage1_regs_3_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_1_4 <= stage1_regs_3_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_1_5 <= stage1_regs_3_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_1_6 <= stage1_regs_3_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_1_7 <= stage1_regs_3_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_3_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_3_1_8 <= stage1_regs_3_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_4_0_0 <= x_n_16; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_0_1 <= stage1_regs_4_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_0_2 <= stage1_regs_4_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_0_3 <= stage1_regs_4_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_0_4 <= stage1_regs_4_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_0_5 <= stage1_regs_4_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_0_6 <= stage1_regs_4_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_0_7 <= stage1_regs_4_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_0_8 <= stage1_regs_4_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_4_1_0 <= a_2_16; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_1_1 <= stage1_regs_4_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_1_2 <= stage1_regs_4_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_1_3 <= stage1_regs_4_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_1_4 <= stage1_regs_4_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_1_5 <= stage1_regs_4_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_1_6 <= stage1_regs_4_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_1_7 <= stage1_regs_4_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_4_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_4_1_8 <= stage1_regs_4_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_5_0_0 <= x_n_20; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_0_1 <= stage1_regs_5_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_0_2 <= stage1_regs_5_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_0_3 <= stage1_regs_5_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_0_4 <= stage1_regs_5_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_0_5 <= stage1_regs_5_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_0_6 <= stage1_regs_5_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_0_7 <= stage1_regs_5_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_0_8 <= stage1_regs_5_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_5_1_0 <= a_2_20; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_1_1 <= stage1_regs_5_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_1_2 <= stage1_regs_5_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_1_3 <= stage1_regs_5_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_1_4 <= stage1_regs_5_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_1_5 <= stage1_regs_5_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_1_6 <= stage1_regs_5_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_1_7 <= stage1_regs_5_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_5_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_5_1_8 <= stage1_regs_5_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_6_0_0 <= x_n_24; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_0_1 <= stage1_regs_6_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_0_2 <= stage1_regs_6_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_0_3 <= stage1_regs_6_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_0_4 <= stage1_regs_6_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_0_5 <= stage1_regs_6_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_0_6 <= stage1_regs_6_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_0_7 <= stage1_regs_6_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_0_8 <= stage1_regs_6_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_6_1_0 <= a_2_24; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_1_1 <= stage1_regs_6_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_1_2 <= stage1_regs_6_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_1_3 <= stage1_regs_6_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_1_4 <= stage1_regs_6_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_1_5 <= stage1_regs_6_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_1_6 <= stage1_regs_6_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_1_7 <= stage1_regs_6_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_6_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_6_1_8 <= stage1_regs_6_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_7_0_0 <= x_n_28; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_0_1 <= stage1_regs_7_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_0_2 <= stage1_regs_7_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_0_3 <= stage1_regs_7_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_0_4 <= stage1_regs_7_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_0_5 <= stage1_regs_7_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_0_6 <= stage1_regs_7_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_0_7 <= stage1_regs_7_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_0_8 <= stage1_regs_7_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_7_1_0 <= a_2_28; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_1_1 <= stage1_regs_7_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_1_2 <= stage1_regs_7_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_1_3 <= stage1_regs_7_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_1_4 <= stage1_regs_7_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_1_5 <= stage1_regs_7_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_1_6 <= stage1_regs_7_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_1_7 <= stage1_regs_7_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_7_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_7_1_8 <= stage1_regs_7_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_8_0_0 <= x_n_32; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_0_1 <= stage1_regs_8_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_0_2 <= stage1_regs_8_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_0_3 <= stage1_regs_8_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_0_4 <= stage1_regs_8_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_0_5 <= stage1_regs_8_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_0_6 <= stage1_regs_8_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_0_7 <= stage1_regs_8_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_0_8 <= stage1_regs_8_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_8_1_0 <= a_2_32; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_1_1 <= stage1_regs_8_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_1_2 <= stage1_regs_8_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_1_3 <= stage1_regs_8_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_1_4 <= stage1_regs_8_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_1_5 <= stage1_regs_8_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_1_6 <= stage1_regs_8_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_1_7 <= stage1_regs_8_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_8_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_8_1_8 <= stage1_regs_8_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_9_0_0 <= x_n_36; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_0_1 <= stage1_regs_9_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_0_2 <= stage1_regs_9_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_0_3 <= stage1_regs_9_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_0_4 <= stage1_regs_9_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_0_5 <= stage1_regs_9_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_0_6 <= stage1_regs_9_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_0_7 <= stage1_regs_9_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_0_8 <= stage1_regs_9_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_9_1_0 <= a_2_36; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_1_1 <= stage1_regs_9_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_1_2 <= stage1_regs_9_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_1_3 <= stage1_regs_9_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_1_4 <= stage1_regs_9_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_1_5 <= stage1_regs_9_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_1_6 <= stage1_regs_9_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_1_7 <= stage1_regs_9_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_9_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_9_1_8 <= stage1_regs_9_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_10_0_0 <= x_n_40; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_0_1 <= stage1_regs_10_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_0_2 <= stage1_regs_10_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_0_3 <= stage1_regs_10_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_0_4 <= stage1_regs_10_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_0_5 <= stage1_regs_10_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_0_6 <= stage1_regs_10_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_0_7 <= stage1_regs_10_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_0_8 <= stage1_regs_10_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_10_1_0 <= a_2_40; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_1_1 <= stage1_regs_10_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_1_2 <= stage1_regs_10_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_1_3 <= stage1_regs_10_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_1_4 <= stage1_regs_10_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_1_5 <= stage1_regs_10_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_1_6 <= stage1_regs_10_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_1_7 <= stage1_regs_10_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_10_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_10_1_8 <= stage1_regs_10_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_11_0_0 <= x_n_44; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_0_1 <= stage1_regs_11_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_0_2 <= stage1_regs_11_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_0_3 <= stage1_regs_11_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_0_4 <= stage1_regs_11_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_0_5 <= stage1_regs_11_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_0_6 <= stage1_regs_11_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_0_7 <= stage1_regs_11_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_0_8 <= stage1_regs_11_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_11_1_0 <= a_2_44; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_1_1 <= stage1_regs_11_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_1_2 <= stage1_regs_11_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_1_3 <= stage1_regs_11_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_1_4 <= stage1_regs_11_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_1_5 <= stage1_regs_11_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_1_6 <= stage1_regs_11_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_1_7 <= stage1_regs_11_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_11_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_11_1_8 <= stage1_regs_11_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_12_0_0 <= x_n_48; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_0_1 <= stage1_regs_12_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_0_2 <= stage1_regs_12_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_0_3 <= stage1_regs_12_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_0_4 <= stage1_regs_12_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_0_5 <= stage1_regs_12_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_0_6 <= stage1_regs_12_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_0_7 <= stage1_regs_12_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_0_8 <= stage1_regs_12_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_12_1_0 <= a_2_48; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_1_1 <= stage1_regs_12_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_1_2 <= stage1_regs_12_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_1_3 <= stage1_regs_12_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_1_4 <= stage1_regs_12_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_1_5 <= stage1_regs_12_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_1_6 <= stage1_regs_12_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_1_7 <= stage1_regs_12_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_12_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_12_1_8 <= stage1_regs_12_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_13_0_0 <= x_n_52; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_0_1 <= stage1_regs_13_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_0_2 <= stage1_regs_13_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_0_3 <= stage1_regs_13_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_0_4 <= stage1_regs_13_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_0_5 <= stage1_regs_13_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_0_6 <= stage1_regs_13_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_0_7 <= stage1_regs_13_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_0_8 <= stage1_regs_13_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_13_1_0 <= a_2_52; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_1_1 <= stage1_regs_13_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_1_2 <= stage1_regs_13_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_1_3 <= stage1_regs_13_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_1_4 <= stage1_regs_13_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_1_5 <= stage1_regs_13_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_1_6 <= stage1_regs_13_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_1_7 <= stage1_regs_13_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_13_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_13_1_8 <= stage1_regs_13_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_14_0_0 <= x_n_56; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_0_1 <= stage1_regs_14_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_0_2 <= stage1_regs_14_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_0_3 <= stage1_regs_14_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_0_4 <= stage1_regs_14_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_0_5 <= stage1_regs_14_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_0_6 <= stage1_regs_14_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_0_7 <= stage1_regs_14_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_0_8 <= stage1_regs_14_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_14_1_0 <= a_2_56; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_1_1 <= stage1_regs_14_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_1_2 <= stage1_regs_14_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_1_3 <= stage1_regs_14_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_1_4 <= stage1_regs_14_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_1_5 <= stage1_regs_14_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_1_6 <= stage1_regs_14_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_1_7 <= stage1_regs_14_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_14_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_14_1_8 <= stage1_regs_14_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_15_0_0 <= x_n_60; // @[FloatingPointDesigns.scala 2018:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_0_1 <= stage1_regs_15_0_0; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_0_2 <= stage1_regs_15_0_1; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_0_3 <= stage1_regs_15_0_2; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_0_4 <= stage1_regs_15_0_3; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_0_5 <= stage1_regs_15_0_4; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_0_6 <= stage1_regs_15_0_5; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_0_7 <= stage1_regs_15_0_6; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_0_8 <= stage1_regs_15_0_7; // @[FloatingPointDesigns.scala 1995:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2015:28]
      stage1_regs_15_1_0 <= a_2_60; // @[FloatingPointDesigns.scala 2019:36]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_1_1 <= stage1_regs_15_1_0; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_1_2 <= stage1_regs_15_1_1; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_1_3 <= stage1_regs_15_1_2; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_1_4 <= stage1_regs_15_1_3; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_1_5 <= stage1_regs_15_1_4; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_1_6 <= stage1_regs_15_1_5; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_1_7 <= stage1_regs_15_1_6; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1980:30]
      stage1_regs_15_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1980:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage1_regs_15_1_8 <= stage1_regs_15_1_7; // @[FloatingPointDesigns.scala 1996:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_0_0_0 <= x_n_1; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_0_1 <= stage2_regs_0_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_0_2 <= stage2_regs_0_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_0_3 <= stage2_regs_0_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_0_4 <= stage2_regs_0_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_0_5 <= stage2_regs_0_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_0_6 <= stage2_regs_0_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_0_7 <= stage2_regs_0_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_0_8 <= stage2_regs_0_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_0_1_0 <= a_2_1; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_1_1 <= stage2_regs_0_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_1_2 <= stage2_regs_0_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_1_3 <= stage2_regs_0_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_1_4 <= stage2_regs_0_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_1_5 <= stage2_regs_0_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_1_6 <= stage2_regs_0_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_1_7 <= stage2_regs_0_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_0_1_8 <= stage2_regs_0_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_1_0_0 <= x_n_5; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_0_1 <= stage2_regs_1_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_0_2 <= stage2_regs_1_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_0_3 <= stage2_regs_1_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_0_4 <= stage2_regs_1_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_0_5 <= stage2_regs_1_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_0_6 <= stage2_regs_1_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_0_7 <= stage2_regs_1_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_0_8 <= stage2_regs_1_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_1_1_0 <= a_2_5; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_1_1 <= stage2_regs_1_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_1_2 <= stage2_regs_1_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_1_3 <= stage2_regs_1_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_1_4 <= stage2_regs_1_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_1_5 <= stage2_regs_1_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_1_6 <= stage2_regs_1_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_1_7 <= stage2_regs_1_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_1_1_8 <= stage2_regs_1_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_2_0_0 <= x_n_9; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_0_1 <= stage2_regs_2_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_0_2 <= stage2_regs_2_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_0_3 <= stage2_regs_2_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_0_4 <= stage2_regs_2_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_0_5 <= stage2_regs_2_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_0_6 <= stage2_regs_2_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_0_7 <= stage2_regs_2_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_0_8 <= stage2_regs_2_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_2_1_0 <= a_2_9; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_1_1 <= stage2_regs_2_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_1_2 <= stage2_regs_2_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_1_3 <= stage2_regs_2_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_1_4 <= stage2_regs_2_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_1_5 <= stage2_regs_2_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_1_6 <= stage2_regs_2_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_1_7 <= stage2_regs_2_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_2_1_8 <= stage2_regs_2_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_3_0_0 <= x_n_13; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_0_1 <= stage2_regs_3_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_0_2 <= stage2_regs_3_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_0_3 <= stage2_regs_3_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_0_4 <= stage2_regs_3_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_0_5 <= stage2_regs_3_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_0_6 <= stage2_regs_3_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_0_7 <= stage2_regs_3_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_0_8 <= stage2_regs_3_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_3_1_0 <= a_2_13; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_1_1 <= stage2_regs_3_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_1_2 <= stage2_regs_3_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_1_3 <= stage2_regs_3_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_1_4 <= stage2_regs_3_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_1_5 <= stage2_regs_3_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_1_6 <= stage2_regs_3_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_1_7 <= stage2_regs_3_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_3_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_3_1_8 <= stage2_regs_3_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_4_0_0 <= x_n_17; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_0_1 <= stage2_regs_4_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_0_2 <= stage2_regs_4_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_0_3 <= stage2_regs_4_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_0_4 <= stage2_regs_4_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_0_5 <= stage2_regs_4_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_0_6 <= stage2_regs_4_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_0_7 <= stage2_regs_4_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_0_8 <= stage2_regs_4_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_4_1_0 <= a_2_17; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_1_1 <= stage2_regs_4_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_1_2 <= stage2_regs_4_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_1_3 <= stage2_regs_4_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_1_4 <= stage2_regs_4_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_1_5 <= stage2_regs_4_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_1_6 <= stage2_regs_4_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_1_7 <= stage2_regs_4_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_4_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_4_1_8 <= stage2_regs_4_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_5_0_0 <= x_n_21; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_0_1 <= stage2_regs_5_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_0_2 <= stage2_regs_5_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_0_3 <= stage2_regs_5_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_0_4 <= stage2_regs_5_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_0_5 <= stage2_regs_5_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_0_6 <= stage2_regs_5_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_0_7 <= stage2_regs_5_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_0_8 <= stage2_regs_5_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_5_1_0 <= a_2_21; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_1_1 <= stage2_regs_5_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_1_2 <= stage2_regs_5_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_1_3 <= stage2_regs_5_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_1_4 <= stage2_regs_5_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_1_5 <= stage2_regs_5_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_1_6 <= stage2_regs_5_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_1_7 <= stage2_regs_5_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_5_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_5_1_8 <= stage2_regs_5_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_6_0_0 <= x_n_25; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_0_1 <= stage2_regs_6_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_0_2 <= stage2_regs_6_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_0_3 <= stage2_regs_6_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_0_4 <= stage2_regs_6_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_0_5 <= stage2_regs_6_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_0_6 <= stage2_regs_6_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_0_7 <= stage2_regs_6_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_0_8 <= stage2_regs_6_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_6_1_0 <= a_2_25; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_1_1 <= stage2_regs_6_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_1_2 <= stage2_regs_6_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_1_3 <= stage2_regs_6_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_1_4 <= stage2_regs_6_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_1_5 <= stage2_regs_6_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_1_6 <= stage2_regs_6_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_1_7 <= stage2_regs_6_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_6_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_6_1_8 <= stage2_regs_6_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_7_0_0 <= x_n_29; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_0_1 <= stage2_regs_7_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_0_2 <= stage2_regs_7_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_0_3 <= stage2_regs_7_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_0_4 <= stage2_regs_7_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_0_5 <= stage2_regs_7_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_0_6 <= stage2_regs_7_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_0_7 <= stage2_regs_7_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_0_8 <= stage2_regs_7_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_7_1_0 <= a_2_29; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_1_1 <= stage2_regs_7_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_1_2 <= stage2_regs_7_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_1_3 <= stage2_regs_7_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_1_4 <= stage2_regs_7_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_1_5 <= stage2_regs_7_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_1_6 <= stage2_regs_7_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_1_7 <= stage2_regs_7_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_7_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_7_1_8 <= stage2_regs_7_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_8_0_0 <= x_n_33; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_0_1 <= stage2_regs_8_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_0_2 <= stage2_regs_8_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_0_3 <= stage2_regs_8_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_0_4 <= stage2_regs_8_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_0_5 <= stage2_regs_8_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_0_6 <= stage2_regs_8_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_0_7 <= stage2_regs_8_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_0_8 <= stage2_regs_8_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_8_1_0 <= a_2_33; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_1_1 <= stage2_regs_8_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_1_2 <= stage2_regs_8_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_1_3 <= stage2_regs_8_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_1_4 <= stage2_regs_8_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_1_5 <= stage2_regs_8_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_1_6 <= stage2_regs_8_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_1_7 <= stage2_regs_8_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_8_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_8_1_8 <= stage2_regs_8_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_9_0_0 <= x_n_37; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_0_1 <= stage2_regs_9_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_0_2 <= stage2_regs_9_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_0_3 <= stage2_regs_9_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_0_4 <= stage2_regs_9_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_0_5 <= stage2_regs_9_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_0_6 <= stage2_regs_9_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_0_7 <= stage2_regs_9_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_0_8 <= stage2_regs_9_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_9_1_0 <= a_2_37; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_1_1 <= stage2_regs_9_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_1_2 <= stage2_regs_9_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_1_3 <= stage2_regs_9_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_1_4 <= stage2_regs_9_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_1_5 <= stage2_regs_9_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_1_6 <= stage2_regs_9_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_1_7 <= stage2_regs_9_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_9_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_9_1_8 <= stage2_regs_9_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_10_0_0 <= x_n_41; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_0_1 <= stage2_regs_10_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_0_2 <= stage2_regs_10_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_0_3 <= stage2_regs_10_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_0_4 <= stage2_regs_10_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_0_5 <= stage2_regs_10_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_0_6 <= stage2_regs_10_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_0_7 <= stage2_regs_10_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_0_8 <= stage2_regs_10_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_10_1_0 <= a_2_41; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_1_1 <= stage2_regs_10_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_1_2 <= stage2_regs_10_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_1_3 <= stage2_regs_10_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_1_4 <= stage2_regs_10_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_1_5 <= stage2_regs_10_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_1_6 <= stage2_regs_10_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_1_7 <= stage2_regs_10_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_10_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_10_1_8 <= stage2_regs_10_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_11_0_0 <= x_n_45; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_0_1 <= stage2_regs_11_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_0_2 <= stage2_regs_11_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_0_3 <= stage2_regs_11_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_0_4 <= stage2_regs_11_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_0_5 <= stage2_regs_11_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_0_6 <= stage2_regs_11_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_0_7 <= stage2_regs_11_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_0_8 <= stage2_regs_11_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_11_1_0 <= a_2_45; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_1_1 <= stage2_regs_11_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_1_2 <= stage2_regs_11_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_1_3 <= stage2_regs_11_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_1_4 <= stage2_regs_11_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_1_5 <= stage2_regs_11_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_1_6 <= stage2_regs_11_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_1_7 <= stage2_regs_11_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_11_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_11_1_8 <= stage2_regs_11_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_12_0_0 <= x_n_49; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_0_1 <= stage2_regs_12_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_0_2 <= stage2_regs_12_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_0_3 <= stage2_regs_12_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_0_4 <= stage2_regs_12_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_0_5 <= stage2_regs_12_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_0_6 <= stage2_regs_12_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_0_7 <= stage2_regs_12_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_0_8 <= stage2_regs_12_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_12_1_0 <= a_2_49; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_1_1 <= stage2_regs_12_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_1_2 <= stage2_regs_12_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_1_3 <= stage2_regs_12_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_1_4 <= stage2_regs_12_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_1_5 <= stage2_regs_12_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_1_6 <= stage2_regs_12_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_1_7 <= stage2_regs_12_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_12_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_12_1_8 <= stage2_regs_12_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_13_0_0 <= x_n_53; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_0_1 <= stage2_regs_13_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_0_2 <= stage2_regs_13_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_0_3 <= stage2_regs_13_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_0_4 <= stage2_regs_13_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_0_5 <= stage2_regs_13_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_0_6 <= stage2_regs_13_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_0_7 <= stage2_regs_13_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_0_8 <= stage2_regs_13_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_13_1_0 <= a_2_53; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_1_1 <= stage2_regs_13_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_1_2 <= stage2_regs_13_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_1_3 <= stage2_regs_13_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_1_4 <= stage2_regs_13_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_1_5 <= stage2_regs_13_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_1_6 <= stage2_regs_13_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_1_7 <= stage2_regs_13_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_13_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_13_1_8 <= stage2_regs_13_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_14_0_0 <= x_n_57; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_0_1 <= stage2_regs_14_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_0_2 <= stage2_regs_14_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_0_3 <= stage2_regs_14_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_0_4 <= stage2_regs_14_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_0_5 <= stage2_regs_14_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_0_6 <= stage2_regs_14_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_0_7 <= stage2_regs_14_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_0_8 <= stage2_regs_14_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_14_1_0 <= a_2_57; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_1_1 <= stage2_regs_14_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_1_2 <= stage2_regs_14_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_1_3 <= stage2_regs_14_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_1_4 <= stage2_regs_14_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_1_5 <= stage2_regs_14_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_1_6 <= stage2_regs_14_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_1_7 <= stage2_regs_14_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_14_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_14_1_8 <= stage2_regs_14_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_15_0_0 <= x_n_61; // @[FloatingPointDesigns.scala 2030:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_0_1 <= stage2_regs_15_0_0; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_0_2 <= stage2_regs_15_0_1; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_0_3 <= stage2_regs_15_0_2; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_0_4 <= stage2_regs_15_0_3; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_0_5 <= stage2_regs_15_0_4; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_0_6 <= stage2_regs_15_0_5; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_0_7 <= stage2_regs_15_0_6; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_0_8 <= stage2_regs_15_0_7; // @[FloatingPointDesigns.scala 1997:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2027:26]
      stage2_regs_15_1_0 <= a_2_61; // @[FloatingPointDesigns.scala 2031:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_1_1 <= stage2_regs_15_1_0; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_1_2 <= stage2_regs_15_1_1; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_1_3 <= stage2_regs_15_1_2; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_1_4 <= stage2_regs_15_1_3; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_1_5 <= stage2_regs_15_1_4; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_1_6 <= stage2_regs_15_1_5; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_1_7 <= stage2_regs_15_1_6; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1981:30]
      stage2_regs_15_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1981:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage2_regs_15_1_8 <= stage2_regs_15_1_7; // @[FloatingPointDesigns.scala 1998:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_0_0_0 <= x_n_2; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_0_1 <= stage3_regs_0_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_0_2 <= stage3_regs_0_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_0_3 <= stage3_regs_0_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_0_4 <= stage3_regs_0_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_0_5 <= stage3_regs_0_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_0_6 <= stage3_regs_0_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_0_7 <= stage3_regs_0_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_0_8 <= stage3_regs_0_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_0_9 <= stage3_regs_0_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_0_10 <= stage3_regs_0_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_0_11 <= stage3_regs_0_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_0_1_0 <= a_2_2; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_1_1 <= stage3_regs_0_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_1_2 <= stage3_regs_0_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_1_3 <= stage3_regs_0_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_1_4 <= stage3_regs_0_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_1_5 <= stage3_regs_0_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_1_6 <= stage3_regs_0_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_1_7 <= stage3_regs_0_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_1_8 <= stage3_regs_0_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_1_9 <= stage3_regs_0_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_1_10 <= stage3_regs_0_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_0_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_0_1_11 <= stage3_regs_0_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_1_0_0 <= x_n_6; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_0_1 <= stage3_regs_1_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_0_2 <= stage3_regs_1_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_0_3 <= stage3_regs_1_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_0_4 <= stage3_regs_1_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_0_5 <= stage3_regs_1_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_0_6 <= stage3_regs_1_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_0_7 <= stage3_regs_1_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_0_8 <= stage3_regs_1_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_0_9 <= stage3_regs_1_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_0_10 <= stage3_regs_1_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_0_11 <= stage3_regs_1_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_1_1_0 <= a_2_6; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_1_1 <= stage3_regs_1_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_1_2 <= stage3_regs_1_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_1_3 <= stage3_regs_1_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_1_4 <= stage3_regs_1_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_1_5 <= stage3_regs_1_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_1_6 <= stage3_regs_1_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_1_7 <= stage3_regs_1_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_1_8 <= stage3_regs_1_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_1_9 <= stage3_regs_1_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_1_10 <= stage3_regs_1_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_1_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_1_1_11 <= stage3_regs_1_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_2_0_0 <= x_n_10; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_0_1 <= stage3_regs_2_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_0_2 <= stage3_regs_2_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_0_3 <= stage3_regs_2_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_0_4 <= stage3_regs_2_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_0_5 <= stage3_regs_2_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_0_6 <= stage3_regs_2_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_0_7 <= stage3_regs_2_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_0_8 <= stage3_regs_2_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_0_9 <= stage3_regs_2_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_0_10 <= stage3_regs_2_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_0_11 <= stage3_regs_2_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_2_1_0 <= a_2_10; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_1_1 <= stage3_regs_2_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_1_2 <= stage3_regs_2_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_1_3 <= stage3_regs_2_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_1_4 <= stage3_regs_2_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_1_5 <= stage3_regs_2_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_1_6 <= stage3_regs_2_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_1_7 <= stage3_regs_2_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_1_8 <= stage3_regs_2_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_1_9 <= stage3_regs_2_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_1_10 <= stage3_regs_2_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_2_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_2_1_11 <= stage3_regs_2_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_3_0_0 <= x_n_14; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_0_1 <= stage3_regs_3_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_0_2 <= stage3_regs_3_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_0_3 <= stage3_regs_3_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_0_4 <= stage3_regs_3_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_0_5 <= stage3_regs_3_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_0_6 <= stage3_regs_3_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_0_7 <= stage3_regs_3_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_0_8 <= stage3_regs_3_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_0_9 <= stage3_regs_3_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_0_10 <= stage3_regs_3_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_0_11 <= stage3_regs_3_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_3_1_0 <= a_2_14; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_1_1 <= stage3_regs_3_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_1_2 <= stage3_regs_3_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_1_3 <= stage3_regs_3_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_1_4 <= stage3_regs_3_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_1_5 <= stage3_regs_3_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_1_6 <= stage3_regs_3_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_1_7 <= stage3_regs_3_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_1_8 <= stage3_regs_3_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_1_9 <= stage3_regs_3_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_1_10 <= stage3_regs_3_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_3_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_3_1_11 <= stage3_regs_3_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_4_0_0 <= x_n_18; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_0_1 <= stage3_regs_4_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_0_2 <= stage3_regs_4_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_0_3 <= stage3_regs_4_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_0_4 <= stage3_regs_4_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_0_5 <= stage3_regs_4_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_0_6 <= stage3_regs_4_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_0_7 <= stage3_regs_4_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_0_8 <= stage3_regs_4_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_0_9 <= stage3_regs_4_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_0_10 <= stage3_regs_4_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_0_11 <= stage3_regs_4_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_4_1_0 <= a_2_18; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_1_1 <= stage3_regs_4_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_1_2 <= stage3_regs_4_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_1_3 <= stage3_regs_4_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_1_4 <= stage3_regs_4_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_1_5 <= stage3_regs_4_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_1_6 <= stage3_regs_4_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_1_7 <= stage3_regs_4_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_1_8 <= stage3_regs_4_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_1_9 <= stage3_regs_4_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_1_10 <= stage3_regs_4_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_4_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_4_1_11 <= stage3_regs_4_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_5_0_0 <= x_n_22; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_0_1 <= stage3_regs_5_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_0_2 <= stage3_regs_5_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_0_3 <= stage3_regs_5_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_0_4 <= stage3_regs_5_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_0_5 <= stage3_regs_5_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_0_6 <= stage3_regs_5_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_0_7 <= stage3_regs_5_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_0_8 <= stage3_regs_5_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_0_9 <= stage3_regs_5_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_0_10 <= stage3_regs_5_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_0_11 <= stage3_regs_5_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_5_1_0 <= a_2_22; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_1_1 <= stage3_regs_5_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_1_2 <= stage3_regs_5_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_1_3 <= stage3_regs_5_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_1_4 <= stage3_regs_5_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_1_5 <= stage3_regs_5_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_1_6 <= stage3_regs_5_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_1_7 <= stage3_regs_5_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_1_8 <= stage3_regs_5_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_1_9 <= stage3_regs_5_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_1_10 <= stage3_regs_5_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_5_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_5_1_11 <= stage3_regs_5_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_6_0_0 <= x_n_26; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_0_1 <= stage3_regs_6_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_0_2 <= stage3_regs_6_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_0_3 <= stage3_regs_6_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_0_4 <= stage3_regs_6_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_0_5 <= stage3_regs_6_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_0_6 <= stage3_regs_6_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_0_7 <= stage3_regs_6_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_0_8 <= stage3_regs_6_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_0_9 <= stage3_regs_6_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_0_10 <= stage3_regs_6_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_0_11 <= stage3_regs_6_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_6_1_0 <= a_2_26; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_1_1 <= stage3_regs_6_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_1_2 <= stage3_regs_6_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_1_3 <= stage3_regs_6_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_1_4 <= stage3_regs_6_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_1_5 <= stage3_regs_6_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_1_6 <= stage3_regs_6_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_1_7 <= stage3_regs_6_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_1_8 <= stage3_regs_6_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_1_9 <= stage3_regs_6_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_1_10 <= stage3_regs_6_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_6_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_6_1_11 <= stage3_regs_6_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_7_0_0 <= x_n_30; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_0_1 <= stage3_regs_7_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_0_2 <= stage3_regs_7_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_0_3 <= stage3_regs_7_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_0_4 <= stage3_regs_7_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_0_5 <= stage3_regs_7_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_0_6 <= stage3_regs_7_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_0_7 <= stage3_regs_7_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_0_8 <= stage3_regs_7_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_0_9 <= stage3_regs_7_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_0_10 <= stage3_regs_7_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_0_11 <= stage3_regs_7_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_7_1_0 <= a_2_30; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_1_1 <= stage3_regs_7_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_1_2 <= stage3_regs_7_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_1_3 <= stage3_regs_7_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_1_4 <= stage3_regs_7_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_1_5 <= stage3_regs_7_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_1_6 <= stage3_regs_7_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_1_7 <= stage3_regs_7_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_1_8 <= stage3_regs_7_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_1_9 <= stage3_regs_7_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_1_10 <= stage3_regs_7_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_7_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_7_1_11 <= stage3_regs_7_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_8_0_0 <= x_n_34; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_0_1 <= stage3_regs_8_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_0_2 <= stage3_regs_8_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_0_3 <= stage3_regs_8_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_0_4 <= stage3_regs_8_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_0_5 <= stage3_regs_8_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_0_6 <= stage3_regs_8_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_0_7 <= stage3_regs_8_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_0_8 <= stage3_regs_8_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_0_9 <= stage3_regs_8_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_0_10 <= stage3_regs_8_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_0_11 <= stage3_regs_8_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_8_1_0 <= a_2_34; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_1_1 <= stage3_regs_8_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_1_2 <= stage3_regs_8_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_1_3 <= stage3_regs_8_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_1_4 <= stage3_regs_8_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_1_5 <= stage3_regs_8_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_1_6 <= stage3_regs_8_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_1_7 <= stage3_regs_8_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_1_8 <= stage3_regs_8_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_1_9 <= stage3_regs_8_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_1_10 <= stage3_regs_8_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_8_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_8_1_11 <= stage3_regs_8_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_9_0_0 <= x_n_38; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_0_1 <= stage3_regs_9_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_0_2 <= stage3_regs_9_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_0_3 <= stage3_regs_9_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_0_4 <= stage3_regs_9_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_0_5 <= stage3_regs_9_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_0_6 <= stage3_regs_9_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_0_7 <= stage3_regs_9_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_0_8 <= stage3_regs_9_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_0_9 <= stage3_regs_9_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_0_10 <= stage3_regs_9_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_0_11 <= stage3_regs_9_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_9_1_0 <= a_2_38; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_1_1 <= stage3_regs_9_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_1_2 <= stage3_regs_9_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_1_3 <= stage3_regs_9_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_1_4 <= stage3_regs_9_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_1_5 <= stage3_regs_9_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_1_6 <= stage3_regs_9_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_1_7 <= stage3_regs_9_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_1_8 <= stage3_regs_9_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_1_9 <= stage3_regs_9_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_1_10 <= stage3_regs_9_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_9_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_9_1_11 <= stage3_regs_9_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_10_0_0 <= x_n_42; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_0_1 <= stage3_regs_10_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_0_2 <= stage3_regs_10_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_0_3 <= stage3_regs_10_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_0_4 <= stage3_regs_10_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_0_5 <= stage3_regs_10_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_0_6 <= stage3_regs_10_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_0_7 <= stage3_regs_10_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_0_8 <= stage3_regs_10_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_0_9 <= stage3_regs_10_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_0_10 <= stage3_regs_10_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_0_11 <= stage3_regs_10_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_10_1_0 <= a_2_42; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_1_1 <= stage3_regs_10_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_1_2 <= stage3_regs_10_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_1_3 <= stage3_regs_10_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_1_4 <= stage3_regs_10_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_1_5 <= stage3_regs_10_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_1_6 <= stage3_regs_10_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_1_7 <= stage3_regs_10_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_1_8 <= stage3_regs_10_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_1_9 <= stage3_regs_10_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_1_10 <= stage3_regs_10_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_10_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_10_1_11 <= stage3_regs_10_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_11_0_0 <= x_n_46; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_0_1 <= stage3_regs_11_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_0_2 <= stage3_regs_11_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_0_3 <= stage3_regs_11_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_0_4 <= stage3_regs_11_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_0_5 <= stage3_regs_11_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_0_6 <= stage3_regs_11_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_0_7 <= stage3_regs_11_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_0_8 <= stage3_regs_11_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_0_9 <= stage3_regs_11_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_0_10 <= stage3_regs_11_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_0_11 <= stage3_regs_11_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_11_1_0 <= a_2_46; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_1_1 <= stage3_regs_11_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_1_2 <= stage3_regs_11_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_1_3 <= stage3_regs_11_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_1_4 <= stage3_regs_11_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_1_5 <= stage3_regs_11_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_1_6 <= stage3_regs_11_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_1_7 <= stage3_regs_11_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_1_8 <= stage3_regs_11_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_1_9 <= stage3_regs_11_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_1_10 <= stage3_regs_11_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_11_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_11_1_11 <= stage3_regs_11_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_12_0_0 <= x_n_50; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_0_1 <= stage3_regs_12_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_0_2 <= stage3_regs_12_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_0_3 <= stage3_regs_12_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_0_4 <= stage3_regs_12_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_0_5 <= stage3_regs_12_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_0_6 <= stage3_regs_12_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_0_7 <= stage3_regs_12_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_0_8 <= stage3_regs_12_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_0_9 <= stage3_regs_12_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_0_10 <= stage3_regs_12_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_0_11 <= stage3_regs_12_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_12_1_0 <= a_2_50; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_1_1 <= stage3_regs_12_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_1_2 <= stage3_regs_12_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_1_3 <= stage3_regs_12_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_1_4 <= stage3_regs_12_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_1_5 <= stage3_regs_12_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_1_6 <= stage3_regs_12_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_1_7 <= stage3_regs_12_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_1_8 <= stage3_regs_12_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_1_9 <= stage3_regs_12_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_1_10 <= stage3_regs_12_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_12_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_12_1_11 <= stage3_regs_12_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_13_0_0 <= x_n_54; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_0_1 <= stage3_regs_13_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_0_2 <= stage3_regs_13_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_0_3 <= stage3_regs_13_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_0_4 <= stage3_regs_13_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_0_5 <= stage3_regs_13_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_0_6 <= stage3_regs_13_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_0_7 <= stage3_regs_13_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_0_8 <= stage3_regs_13_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_0_9 <= stage3_regs_13_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_0_10 <= stage3_regs_13_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_0_11 <= stage3_regs_13_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_13_1_0 <= a_2_54; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_1_1 <= stage3_regs_13_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_1_2 <= stage3_regs_13_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_1_3 <= stage3_regs_13_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_1_4 <= stage3_regs_13_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_1_5 <= stage3_regs_13_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_1_6 <= stage3_regs_13_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_1_7 <= stage3_regs_13_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_1_8 <= stage3_regs_13_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_1_9 <= stage3_regs_13_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_1_10 <= stage3_regs_13_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_13_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_13_1_11 <= stage3_regs_13_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_14_0_0 <= x_n_58; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_0_1 <= stage3_regs_14_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_0_2 <= stage3_regs_14_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_0_3 <= stage3_regs_14_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_0_4 <= stage3_regs_14_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_0_5 <= stage3_regs_14_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_0_6 <= stage3_regs_14_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_0_7 <= stage3_regs_14_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_0_8 <= stage3_regs_14_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_0_9 <= stage3_regs_14_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_0_10 <= stage3_regs_14_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_0_11 <= stage3_regs_14_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_14_1_0 <= a_2_58; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_1_1 <= stage3_regs_14_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_1_2 <= stage3_regs_14_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_1_3 <= stage3_regs_14_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_1_4 <= stage3_regs_14_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_1_5 <= stage3_regs_14_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_1_6 <= stage3_regs_14_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_1_7 <= stage3_regs_14_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_1_8 <= stage3_regs_14_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_1_9 <= stage3_regs_14_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_1_10 <= stage3_regs_14_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_14_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_14_1_11 <= stage3_regs_14_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_15_0_0 <= x_n_62; // @[FloatingPointDesigns.scala 2039:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_0_1 <= stage3_regs_15_0_0; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_0_2 <= stage3_regs_15_0_1; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_0_3 <= stage3_regs_15_0_2; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_0_4 <= stage3_regs_15_0_3; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_0_5 <= stage3_regs_15_0_4; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_0_6 <= stage3_regs_15_0_5; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_0_7 <= stage3_regs_15_0_6; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_0_8 <= stage3_regs_15_0_7; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_0_9 <= stage3_regs_15_0_8; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_0_10 <= stage3_regs_15_0_9; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_0_11 <= stage3_regs_15_0_10; // @[FloatingPointDesigns.scala 1992:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2036:26]
      stage3_regs_15_1_0 <= a_2_62; // @[FloatingPointDesigns.scala 2040:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_1_1 <= stage3_regs_15_1_0; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_1_2 <= stage3_regs_15_1_1; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_1_3 <= stage3_regs_15_1_2; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_1_4 <= stage3_regs_15_1_3; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_1_5 <= stage3_regs_15_1_4; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_1_6 <= stage3_regs_15_1_5; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_1_7 <= stage3_regs_15_1_6; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_1_8 <= stage3_regs_15_1_7; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_1_9 <= stage3_regs_15_1_8; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_1_10 <= stage3_regs_15_1_9; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1982:30]
      stage3_regs_15_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1982:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage3_regs_15_1_11 <= stage3_regs_15_1_10; // @[FloatingPointDesigns.scala 1993:32]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_0_1_0 <= a_2_3; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_0_1_1 <= stage4_regs_0_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_0_1_2 <= stage4_regs_0_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_0_1_3 <= stage4_regs_0_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_0_1_4 <= stage4_regs_0_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_0_1_5 <= stage4_regs_0_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_0_1_6 <= stage4_regs_0_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_0_1_7 <= stage4_regs_0_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_0_1_8 <= stage4_regs_0_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_1_1_0 <= a_2_7; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_1_1_1 <= stage4_regs_1_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_1_1_2 <= stage4_regs_1_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_1_1_3 <= stage4_regs_1_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_1_1_4 <= stage4_regs_1_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_1_1_5 <= stage4_regs_1_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_1_1_6 <= stage4_regs_1_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_1_1_7 <= stage4_regs_1_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_1_1_8 <= stage4_regs_1_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_2_1_0 <= a_2_11; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_2_1_1 <= stage4_regs_2_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_2_1_2 <= stage4_regs_2_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_2_1_3 <= stage4_regs_2_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_2_1_4 <= stage4_regs_2_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_2_1_5 <= stage4_regs_2_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_2_1_6 <= stage4_regs_2_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_2_1_7 <= stage4_regs_2_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_2_1_8 <= stage4_regs_2_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_3_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_3_1_0 <= a_2_15; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_3_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_3_1_1 <= stage4_regs_3_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_3_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_3_1_2 <= stage4_regs_3_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_3_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_3_1_3 <= stage4_regs_3_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_3_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_3_1_4 <= stage4_regs_3_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_3_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_3_1_5 <= stage4_regs_3_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_3_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_3_1_6 <= stage4_regs_3_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_3_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_3_1_7 <= stage4_regs_3_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_3_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_3_1_8 <= stage4_regs_3_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_4_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_4_1_0 <= a_2_19; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_4_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_4_1_1 <= stage4_regs_4_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_4_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_4_1_2 <= stage4_regs_4_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_4_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_4_1_3 <= stage4_regs_4_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_4_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_4_1_4 <= stage4_regs_4_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_4_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_4_1_5 <= stage4_regs_4_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_4_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_4_1_6 <= stage4_regs_4_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_4_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_4_1_7 <= stage4_regs_4_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_4_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_4_1_8 <= stage4_regs_4_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_5_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_5_1_0 <= a_2_23; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_5_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_5_1_1 <= stage4_regs_5_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_5_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_5_1_2 <= stage4_regs_5_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_5_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_5_1_3 <= stage4_regs_5_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_5_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_5_1_4 <= stage4_regs_5_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_5_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_5_1_5 <= stage4_regs_5_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_5_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_5_1_6 <= stage4_regs_5_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_5_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_5_1_7 <= stage4_regs_5_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_5_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_5_1_8 <= stage4_regs_5_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_6_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_6_1_0 <= a_2_27; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_6_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_6_1_1 <= stage4_regs_6_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_6_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_6_1_2 <= stage4_regs_6_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_6_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_6_1_3 <= stage4_regs_6_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_6_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_6_1_4 <= stage4_regs_6_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_6_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_6_1_5 <= stage4_regs_6_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_6_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_6_1_6 <= stage4_regs_6_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_6_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_6_1_7 <= stage4_regs_6_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_6_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_6_1_8 <= stage4_regs_6_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_7_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_7_1_0 <= a_2_31; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_7_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_7_1_1 <= stage4_regs_7_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_7_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_7_1_2 <= stage4_regs_7_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_7_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_7_1_3 <= stage4_regs_7_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_7_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_7_1_4 <= stage4_regs_7_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_7_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_7_1_5 <= stage4_regs_7_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_7_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_7_1_6 <= stage4_regs_7_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_7_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_7_1_7 <= stage4_regs_7_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_7_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_7_1_8 <= stage4_regs_7_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_8_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_8_1_0 <= a_2_35; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_8_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_8_1_1 <= stage4_regs_8_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_8_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_8_1_2 <= stage4_regs_8_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_8_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_8_1_3 <= stage4_regs_8_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_8_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_8_1_4 <= stage4_regs_8_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_8_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_8_1_5 <= stage4_regs_8_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_8_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_8_1_6 <= stage4_regs_8_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_8_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_8_1_7 <= stage4_regs_8_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_8_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_8_1_8 <= stage4_regs_8_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_9_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_9_1_0 <= a_2_39; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_9_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_9_1_1 <= stage4_regs_9_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_9_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_9_1_2 <= stage4_regs_9_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_9_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_9_1_3 <= stage4_regs_9_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_9_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_9_1_4 <= stage4_regs_9_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_9_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_9_1_5 <= stage4_regs_9_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_9_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_9_1_6 <= stage4_regs_9_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_9_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_9_1_7 <= stage4_regs_9_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_9_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_9_1_8 <= stage4_regs_9_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_10_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_10_1_0 <= a_2_43; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_10_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_10_1_1 <= stage4_regs_10_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_10_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_10_1_2 <= stage4_regs_10_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_10_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_10_1_3 <= stage4_regs_10_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_10_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_10_1_4 <= stage4_regs_10_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_10_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_10_1_5 <= stage4_regs_10_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_10_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_10_1_6 <= stage4_regs_10_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_10_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_10_1_7 <= stage4_regs_10_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_10_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_10_1_8 <= stage4_regs_10_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_11_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_11_1_0 <= a_2_47; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_11_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_11_1_1 <= stage4_regs_11_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_11_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_11_1_2 <= stage4_regs_11_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_11_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_11_1_3 <= stage4_regs_11_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_11_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_11_1_4 <= stage4_regs_11_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_11_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_11_1_5 <= stage4_regs_11_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_11_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_11_1_6 <= stage4_regs_11_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_11_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_11_1_7 <= stage4_regs_11_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_11_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_11_1_8 <= stage4_regs_11_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_12_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_12_1_0 <= a_2_51; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_12_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_12_1_1 <= stage4_regs_12_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_12_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_12_1_2 <= stage4_regs_12_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_12_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_12_1_3 <= stage4_regs_12_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_12_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_12_1_4 <= stage4_regs_12_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_12_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_12_1_5 <= stage4_regs_12_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_12_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_12_1_6 <= stage4_regs_12_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_12_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_12_1_7 <= stage4_regs_12_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_12_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_12_1_8 <= stage4_regs_12_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_13_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_13_1_0 <= a_2_55; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_13_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_13_1_1 <= stage4_regs_13_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_13_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_13_1_2 <= stage4_regs_13_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_13_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_13_1_3 <= stage4_regs_13_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_13_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_13_1_4 <= stage4_regs_13_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_13_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_13_1_5 <= stage4_regs_13_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_13_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_13_1_6 <= stage4_regs_13_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_13_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_13_1_7 <= stage4_regs_13_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_13_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_13_1_8 <= stage4_regs_13_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_14_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_14_1_0 <= a_2_59; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_14_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_14_1_1 <= stage4_regs_14_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_14_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_14_1_2 <= stage4_regs_14_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_14_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_14_1_3 <= stage4_regs_14_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_14_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_14_1_4 <= stage4_regs_14_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_14_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_14_1_5 <= stage4_regs_14_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_14_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_14_1_6 <= stage4_regs_14_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_14_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_14_1_7 <= stage4_regs_14_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_14_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_14_1_8 <= stage4_regs_14_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_15_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 2045:26]
      stage4_regs_15_1_0 <= a_2_63; // @[FloatingPointDesigns.scala 2047:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_15_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_15_1_1 <= stage4_regs_15_1_0; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_15_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_15_1_2 <= stage4_regs_15_1_1; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_15_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_15_1_3 <= stage4_regs_15_1_2; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_15_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_15_1_4 <= stage4_regs_15_1_3; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_15_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_15_1_5 <= stage4_regs_15_1_4; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_15_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_15_1_6 <= stage4_regs_15_1_5; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_15_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_15_1_7 <= stage4_regs_15_1_6; // @[FloatingPointDesigns.scala 1999:34]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1983:30]
      stage4_regs_15_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1983:30]
    end else if (io_in_en) begin // @[FloatingPointDesigns.scala 1990:22]
      stage4_regs_15_1_8 <= stage4_regs_15_1_7; // @[FloatingPointDesigns.scala 1999:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  x_n_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  x_n_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  x_n_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  x_n_4 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  x_n_5 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  x_n_6 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  x_n_8 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  x_n_9 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  x_n_10 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  x_n_12 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  x_n_13 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  x_n_14 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  x_n_16 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  x_n_17 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  x_n_18 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  x_n_20 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  x_n_21 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  x_n_22 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  x_n_24 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  x_n_25 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  x_n_26 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  x_n_28 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  x_n_29 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  x_n_30 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  x_n_32 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  x_n_33 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  x_n_34 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  x_n_36 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  x_n_37 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  x_n_38 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  x_n_40 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  x_n_41 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  x_n_42 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  x_n_44 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  x_n_45 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  x_n_46 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  x_n_48 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  x_n_49 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  x_n_50 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  x_n_52 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  x_n_53 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  x_n_54 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  x_n_56 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  x_n_57 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  x_n_58 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  x_n_60 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  x_n_61 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  x_n_62 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  a_2_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  a_2_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  a_2_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  a_2_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  a_2_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  a_2_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  a_2_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  a_2_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  a_2_8 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  a_2_9 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  a_2_10 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  a_2_11 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  a_2_12 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  a_2_13 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  a_2_14 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  a_2_15 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  a_2_16 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  a_2_17 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  a_2_18 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  a_2_19 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  a_2_20 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  a_2_21 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  a_2_22 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  a_2_23 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  a_2_24 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  a_2_25 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  a_2_26 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  a_2_27 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  a_2_28 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  a_2_29 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  a_2_30 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  a_2_31 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  a_2_32 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  a_2_33 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  a_2_34 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  a_2_35 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  a_2_36 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  a_2_37 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  a_2_38 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  a_2_39 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  a_2_40 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  a_2_41 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  a_2_42 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  a_2_43 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  a_2_44 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  a_2_45 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  a_2_46 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  a_2_47 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  a_2_48 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  a_2_49 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  a_2_50 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  a_2_51 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  a_2_52 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  a_2_53 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  a_2_54 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  a_2_55 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  a_2_56 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  a_2_57 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  a_2_58 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  a_2_59 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  a_2_60 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  a_2_61 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  a_2_62 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  a_2_63 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  stage1_regs_0_0_0 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  stage1_regs_0_0_1 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  stage1_regs_0_0_2 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  stage1_regs_0_0_3 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  stage1_regs_0_0_4 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  stage1_regs_0_0_5 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  stage1_regs_0_0_6 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  stage1_regs_0_0_7 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  stage1_regs_0_0_8 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  stage1_regs_0_1_0 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  stage1_regs_0_1_1 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  stage1_regs_0_1_2 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  stage1_regs_0_1_3 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  stage1_regs_0_1_4 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  stage1_regs_0_1_5 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  stage1_regs_0_1_6 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  stage1_regs_0_1_7 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  stage1_regs_0_1_8 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  stage1_regs_1_0_0 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  stage1_regs_1_0_1 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  stage1_regs_1_0_2 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  stage1_regs_1_0_3 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  stage1_regs_1_0_4 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  stage1_regs_1_0_5 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  stage1_regs_1_0_6 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  stage1_regs_1_0_7 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  stage1_regs_1_0_8 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  stage1_regs_1_1_0 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  stage1_regs_1_1_1 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  stage1_regs_1_1_2 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  stage1_regs_1_1_3 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  stage1_regs_1_1_4 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  stage1_regs_1_1_5 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  stage1_regs_1_1_6 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  stage1_regs_1_1_7 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  stage1_regs_1_1_8 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  stage1_regs_2_0_0 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  stage1_regs_2_0_1 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  stage1_regs_2_0_2 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  stage1_regs_2_0_3 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  stage1_regs_2_0_4 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  stage1_regs_2_0_5 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  stage1_regs_2_0_6 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  stage1_regs_2_0_7 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  stage1_regs_2_0_8 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  stage1_regs_2_1_0 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  stage1_regs_2_1_1 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  stage1_regs_2_1_2 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  stage1_regs_2_1_3 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  stage1_regs_2_1_4 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  stage1_regs_2_1_5 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  stage1_regs_2_1_6 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  stage1_regs_2_1_7 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  stage1_regs_2_1_8 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  stage1_regs_3_0_0 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  stage1_regs_3_0_1 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  stage1_regs_3_0_2 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  stage1_regs_3_0_3 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  stage1_regs_3_0_4 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  stage1_regs_3_0_5 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  stage1_regs_3_0_6 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  stage1_regs_3_0_7 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  stage1_regs_3_0_8 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  stage1_regs_3_1_0 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  stage1_regs_3_1_1 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  stage1_regs_3_1_2 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  stage1_regs_3_1_3 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  stage1_regs_3_1_4 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  stage1_regs_3_1_5 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  stage1_regs_3_1_6 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  stage1_regs_3_1_7 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  stage1_regs_3_1_8 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  stage1_regs_4_0_0 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  stage1_regs_4_0_1 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  stage1_regs_4_0_2 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  stage1_regs_4_0_3 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  stage1_regs_4_0_4 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  stage1_regs_4_0_5 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  stage1_regs_4_0_6 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  stage1_regs_4_0_7 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  stage1_regs_4_0_8 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  stage1_regs_4_1_0 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  stage1_regs_4_1_1 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  stage1_regs_4_1_2 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  stage1_regs_4_1_3 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  stage1_regs_4_1_4 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  stage1_regs_4_1_5 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  stage1_regs_4_1_6 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  stage1_regs_4_1_7 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  stage1_regs_4_1_8 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  stage1_regs_5_0_0 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  stage1_regs_5_0_1 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  stage1_regs_5_0_2 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  stage1_regs_5_0_3 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  stage1_regs_5_0_4 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  stage1_regs_5_0_5 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  stage1_regs_5_0_6 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  stage1_regs_5_0_7 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  stage1_regs_5_0_8 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  stage1_regs_5_1_0 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  stage1_regs_5_1_1 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  stage1_regs_5_1_2 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  stage1_regs_5_1_3 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  stage1_regs_5_1_4 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  stage1_regs_5_1_5 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  stage1_regs_5_1_6 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  stage1_regs_5_1_7 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  stage1_regs_5_1_8 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  stage1_regs_6_0_0 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  stage1_regs_6_0_1 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  stage1_regs_6_0_2 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  stage1_regs_6_0_3 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  stage1_regs_6_0_4 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  stage1_regs_6_0_5 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  stage1_regs_6_0_6 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  stage1_regs_6_0_7 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  stage1_regs_6_0_8 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  stage1_regs_6_1_0 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  stage1_regs_6_1_1 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  stage1_regs_6_1_2 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  stage1_regs_6_1_3 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  stage1_regs_6_1_4 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  stage1_regs_6_1_5 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  stage1_regs_6_1_6 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  stage1_regs_6_1_7 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  stage1_regs_6_1_8 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  stage1_regs_7_0_0 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  stage1_regs_7_0_1 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  stage1_regs_7_0_2 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  stage1_regs_7_0_3 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  stage1_regs_7_0_4 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  stage1_regs_7_0_5 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  stage1_regs_7_0_6 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  stage1_regs_7_0_7 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  stage1_regs_7_0_8 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  stage1_regs_7_1_0 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  stage1_regs_7_1_1 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  stage1_regs_7_1_2 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  stage1_regs_7_1_3 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  stage1_regs_7_1_4 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  stage1_regs_7_1_5 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  stage1_regs_7_1_6 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  stage1_regs_7_1_7 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  stage1_regs_7_1_8 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  stage1_regs_8_0_0 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  stage1_regs_8_0_1 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  stage1_regs_8_0_2 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  stage1_regs_8_0_3 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  stage1_regs_8_0_4 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  stage1_regs_8_0_5 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  stage1_regs_8_0_6 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  stage1_regs_8_0_7 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  stage1_regs_8_0_8 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  stage1_regs_8_1_0 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  stage1_regs_8_1_1 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  stage1_regs_8_1_2 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  stage1_regs_8_1_3 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  stage1_regs_8_1_4 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  stage1_regs_8_1_5 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  stage1_regs_8_1_6 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  stage1_regs_8_1_7 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  stage1_regs_8_1_8 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  stage1_regs_9_0_0 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  stage1_regs_9_0_1 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  stage1_regs_9_0_2 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  stage1_regs_9_0_3 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  stage1_regs_9_0_4 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  stage1_regs_9_0_5 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  stage1_regs_9_0_6 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  stage1_regs_9_0_7 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  stage1_regs_9_0_8 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  stage1_regs_9_1_0 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  stage1_regs_9_1_1 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  stage1_regs_9_1_2 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  stage1_regs_9_1_3 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  stage1_regs_9_1_4 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  stage1_regs_9_1_5 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  stage1_regs_9_1_6 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  stage1_regs_9_1_7 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  stage1_regs_9_1_8 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  stage1_regs_10_0_0 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  stage1_regs_10_0_1 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  stage1_regs_10_0_2 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  stage1_regs_10_0_3 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  stage1_regs_10_0_4 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  stage1_regs_10_0_5 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  stage1_regs_10_0_6 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  stage1_regs_10_0_7 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  stage1_regs_10_0_8 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  stage1_regs_10_1_0 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  stage1_regs_10_1_1 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  stage1_regs_10_1_2 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  stage1_regs_10_1_3 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  stage1_regs_10_1_4 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  stage1_regs_10_1_5 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  stage1_regs_10_1_6 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  stage1_regs_10_1_7 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  stage1_regs_10_1_8 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  stage1_regs_11_0_0 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  stage1_regs_11_0_1 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  stage1_regs_11_0_2 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  stage1_regs_11_0_3 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  stage1_regs_11_0_4 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  stage1_regs_11_0_5 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  stage1_regs_11_0_6 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  stage1_regs_11_0_7 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  stage1_regs_11_0_8 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  stage1_regs_11_1_0 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  stage1_regs_11_1_1 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  stage1_regs_11_1_2 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  stage1_regs_11_1_3 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  stage1_regs_11_1_4 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  stage1_regs_11_1_5 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  stage1_regs_11_1_6 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  stage1_regs_11_1_7 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  stage1_regs_11_1_8 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  stage1_regs_12_0_0 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  stage1_regs_12_0_1 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  stage1_regs_12_0_2 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  stage1_regs_12_0_3 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  stage1_regs_12_0_4 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  stage1_regs_12_0_5 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  stage1_regs_12_0_6 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  stage1_regs_12_0_7 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  stage1_regs_12_0_8 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  stage1_regs_12_1_0 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  stage1_regs_12_1_1 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  stage1_regs_12_1_2 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  stage1_regs_12_1_3 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  stage1_regs_12_1_4 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  stage1_regs_12_1_5 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  stage1_regs_12_1_6 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  stage1_regs_12_1_7 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  stage1_regs_12_1_8 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  stage1_regs_13_0_0 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  stage1_regs_13_0_1 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  stage1_regs_13_0_2 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  stage1_regs_13_0_3 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  stage1_regs_13_0_4 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  stage1_regs_13_0_5 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  stage1_regs_13_0_6 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  stage1_regs_13_0_7 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  stage1_regs_13_0_8 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  stage1_regs_13_1_0 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  stage1_regs_13_1_1 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  stage1_regs_13_1_2 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  stage1_regs_13_1_3 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  stage1_regs_13_1_4 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  stage1_regs_13_1_5 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  stage1_regs_13_1_6 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  stage1_regs_13_1_7 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  stage1_regs_13_1_8 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  stage1_regs_14_0_0 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  stage1_regs_14_0_1 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  stage1_regs_14_0_2 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  stage1_regs_14_0_3 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  stage1_regs_14_0_4 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  stage1_regs_14_0_5 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  stage1_regs_14_0_6 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  stage1_regs_14_0_7 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  stage1_regs_14_0_8 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  stage1_regs_14_1_0 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  stage1_regs_14_1_1 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  stage1_regs_14_1_2 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  stage1_regs_14_1_3 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  stage1_regs_14_1_4 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  stage1_regs_14_1_5 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  stage1_regs_14_1_6 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  stage1_regs_14_1_7 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  stage1_regs_14_1_8 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  stage1_regs_15_0_0 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  stage1_regs_15_0_1 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  stage1_regs_15_0_2 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  stage1_regs_15_0_3 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  stage1_regs_15_0_4 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  stage1_regs_15_0_5 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  stage1_regs_15_0_6 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  stage1_regs_15_0_7 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  stage1_regs_15_0_8 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  stage1_regs_15_1_0 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  stage1_regs_15_1_1 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  stage1_regs_15_1_2 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  stage1_regs_15_1_3 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  stage1_regs_15_1_4 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  stage1_regs_15_1_5 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  stage1_regs_15_1_6 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  stage1_regs_15_1_7 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  stage1_regs_15_1_8 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  stage2_regs_0_0_0 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  stage2_regs_0_0_1 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  stage2_regs_0_0_2 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  stage2_regs_0_0_3 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  stage2_regs_0_0_4 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  stage2_regs_0_0_5 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  stage2_regs_0_0_6 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  stage2_regs_0_0_7 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  stage2_regs_0_0_8 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  stage2_regs_0_1_0 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  stage2_regs_0_1_1 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  stage2_regs_0_1_2 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  stage2_regs_0_1_3 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  stage2_regs_0_1_4 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  stage2_regs_0_1_5 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  stage2_regs_0_1_6 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  stage2_regs_0_1_7 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  stage2_regs_0_1_8 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  stage2_regs_1_0_0 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  stage2_regs_1_0_1 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  stage2_regs_1_0_2 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  stage2_regs_1_0_3 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  stage2_regs_1_0_4 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  stage2_regs_1_0_5 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  stage2_regs_1_0_6 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  stage2_regs_1_0_7 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  stage2_regs_1_0_8 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  stage2_regs_1_1_0 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  stage2_regs_1_1_1 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  stage2_regs_1_1_2 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  stage2_regs_1_1_3 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  stage2_regs_1_1_4 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  stage2_regs_1_1_5 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  stage2_regs_1_1_6 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  stage2_regs_1_1_7 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  stage2_regs_1_1_8 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  stage2_regs_2_0_0 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  stage2_regs_2_0_1 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  stage2_regs_2_0_2 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  stage2_regs_2_0_3 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  stage2_regs_2_0_4 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  stage2_regs_2_0_5 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  stage2_regs_2_0_6 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  stage2_regs_2_0_7 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  stage2_regs_2_0_8 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  stage2_regs_2_1_0 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  stage2_regs_2_1_1 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  stage2_regs_2_1_2 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  stage2_regs_2_1_3 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  stage2_regs_2_1_4 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  stage2_regs_2_1_5 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  stage2_regs_2_1_6 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  stage2_regs_2_1_7 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  stage2_regs_2_1_8 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  stage2_regs_3_0_0 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  stage2_regs_3_0_1 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  stage2_regs_3_0_2 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  stage2_regs_3_0_3 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  stage2_regs_3_0_4 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  stage2_regs_3_0_5 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  stage2_regs_3_0_6 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  stage2_regs_3_0_7 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  stage2_regs_3_0_8 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  stage2_regs_3_1_0 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  stage2_regs_3_1_1 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  stage2_regs_3_1_2 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  stage2_regs_3_1_3 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  stage2_regs_3_1_4 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  stage2_regs_3_1_5 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  stage2_regs_3_1_6 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  stage2_regs_3_1_7 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  stage2_regs_3_1_8 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  stage2_regs_4_0_0 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  stage2_regs_4_0_1 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  stage2_regs_4_0_2 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  stage2_regs_4_0_3 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  stage2_regs_4_0_4 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  stage2_regs_4_0_5 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  stage2_regs_4_0_6 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  stage2_regs_4_0_7 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  stage2_regs_4_0_8 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  stage2_regs_4_1_0 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  stage2_regs_4_1_1 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  stage2_regs_4_1_2 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  stage2_regs_4_1_3 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  stage2_regs_4_1_4 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  stage2_regs_4_1_5 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  stage2_regs_4_1_6 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  stage2_regs_4_1_7 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  stage2_regs_4_1_8 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  stage2_regs_5_0_0 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  stage2_regs_5_0_1 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  stage2_regs_5_0_2 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  stage2_regs_5_0_3 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  stage2_regs_5_0_4 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  stage2_regs_5_0_5 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  stage2_regs_5_0_6 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  stage2_regs_5_0_7 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  stage2_regs_5_0_8 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  stage2_regs_5_1_0 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  stage2_regs_5_1_1 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  stage2_regs_5_1_2 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  stage2_regs_5_1_3 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  stage2_regs_5_1_4 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  stage2_regs_5_1_5 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  stage2_regs_5_1_6 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  stage2_regs_5_1_7 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  stage2_regs_5_1_8 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  stage2_regs_6_0_0 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  stage2_regs_6_0_1 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  stage2_regs_6_0_2 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  stage2_regs_6_0_3 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  stage2_regs_6_0_4 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  stage2_regs_6_0_5 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  stage2_regs_6_0_6 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  stage2_regs_6_0_7 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  stage2_regs_6_0_8 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  stage2_regs_6_1_0 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  stage2_regs_6_1_1 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  stage2_regs_6_1_2 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  stage2_regs_6_1_3 = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  stage2_regs_6_1_4 = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  stage2_regs_6_1_5 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  stage2_regs_6_1_6 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  stage2_regs_6_1_7 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  stage2_regs_6_1_8 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  stage2_regs_7_0_0 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  stage2_regs_7_0_1 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  stage2_regs_7_0_2 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  stage2_regs_7_0_3 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  stage2_regs_7_0_4 = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  stage2_regs_7_0_5 = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  stage2_regs_7_0_6 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  stage2_regs_7_0_7 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  stage2_regs_7_0_8 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  stage2_regs_7_1_0 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  stage2_regs_7_1_1 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  stage2_regs_7_1_2 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  stage2_regs_7_1_3 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  stage2_regs_7_1_4 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  stage2_regs_7_1_5 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  stage2_regs_7_1_6 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  stage2_regs_7_1_7 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  stage2_regs_7_1_8 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  stage2_regs_8_0_0 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  stage2_regs_8_0_1 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  stage2_regs_8_0_2 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  stage2_regs_8_0_3 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  stage2_regs_8_0_4 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  stage2_regs_8_0_5 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  stage2_regs_8_0_6 = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  stage2_regs_8_0_7 = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  stage2_regs_8_0_8 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  stage2_regs_8_1_0 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  stage2_regs_8_1_1 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  stage2_regs_8_1_2 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  stage2_regs_8_1_3 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  stage2_regs_8_1_4 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  stage2_regs_8_1_5 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  stage2_regs_8_1_6 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  stage2_regs_8_1_7 = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  stage2_regs_8_1_8 = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  stage2_regs_9_0_0 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  stage2_regs_9_0_1 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  stage2_regs_9_0_2 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  stage2_regs_9_0_3 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  stage2_regs_9_0_4 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  stage2_regs_9_0_5 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  stage2_regs_9_0_6 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  stage2_regs_9_0_7 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  stage2_regs_9_0_8 = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  stage2_regs_9_1_0 = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  stage2_regs_9_1_1 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  stage2_regs_9_1_2 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  stage2_regs_9_1_3 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  stage2_regs_9_1_4 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  stage2_regs_9_1_5 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  stage2_regs_9_1_6 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  stage2_regs_9_1_7 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  stage2_regs_9_1_8 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  stage2_regs_10_0_0 = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  stage2_regs_10_0_1 = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  stage2_regs_10_0_2 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  stage2_regs_10_0_3 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  stage2_regs_10_0_4 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  stage2_regs_10_0_5 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  stage2_regs_10_0_6 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  stage2_regs_10_0_7 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  stage2_regs_10_0_8 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  stage2_regs_10_1_0 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  stage2_regs_10_1_1 = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  stage2_regs_10_1_2 = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  stage2_regs_10_1_3 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  stage2_regs_10_1_4 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  stage2_regs_10_1_5 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  stage2_regs_10_1_6 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  stage2_regs_10_1_7 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  stage2_regs_10_1_8 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  stage2_regs_11_0_0 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  stage2_regs_11_0_1 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  stage2_regs_11_0_2 = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  stage2_regs_11_0_3 = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  stage2_regs_11_0_4 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  stage2_regs_11_0_5 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  stage2_regs_11_0_6 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  stage2_regs_11_0_7 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  stage2_regs_11_0_8 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  stage2_regs_11_1_0 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  stage2_regs_11_1_1 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  stage2_regs_11_1_2 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  stage2_regs_11_1_3 = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  stage2_regs_11_1_4 = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  stage2_regs_11_1_5 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  stage2_regs_11_1_6 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  stage2_regs_11_1_7 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  stage2_regs_11_1_8 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  stage2_regs_12_0_0 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  stage2_regs_12_0_1 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  stage2_regs_12_0_2 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  stage2_regs_12_0_3 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  stage2_regs_12_0_4 = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  stage2_regs_12_0_5 = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  stage2_regs_12_0_6 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  stage2_regs_12_0_7 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  stage2_regs_12_0_8 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  stage2_regs_12_1_0 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  stage2_regs_12_1_1 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  stage2_regs_12_1_2 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  stage2_regs_12_1_3 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  stage2_regs_12_1_4 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  stage2_regs_12_1_5 = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  stage2_regs_12_1_6 = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  stage2_regs_12_1_7 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  stage2_regs_12_1_8 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  stage2_regs_13_0_0 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  stage2_regs_13_0_1 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  stage2_regs_13_0_2 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  stage2_regs_13_0_3 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  stage2_regs_13_0_4 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  stage2_regs_13_0_5 = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  stage2_regs_13_0_6 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  stage2_regs_13_0_7 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  stage2_regs_13_0_8 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  stage2_regs_13_1_0 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  stage2_regs_13_1_1 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  stage2_regs_13_1_2 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  stage2_regs_13_1_3 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  stage2_regs_13_1_4 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  stage2_regs_13_1_5 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  stage2_regs_13_1_6 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  stage2_regs_13_1_7 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  stage2_regs_13_1_8 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  stage2_regs_14_0_0 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  stage2_regs_14_0_1 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  stage2_regs_14_0_2 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  stage2_regs_14_0_3 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  stage2_regs_14_0_4 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  stage2_regs_14_0_5 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  stage2_regs_14_0_6 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  stage2_regs_14_0_7 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  stage2_regs_14_0_8 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  stage2_regs_14_1_0 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  stage2_regs_14_1_1 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  stage2_regs_14_1_2 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  stage2_regs_14_1_3 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  stage2_regs_14_1_4 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  stage2_regs_14_1_5 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  stage2_regs_14_1_6 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  stage2_regs_14_1_7 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  stage2_regs_14_1_8 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  stage2_regs_15_0_0 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  stage2_regs_15_0_1 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  stage2_regs_15_0_2 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  stage2_regs_15_0_3 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  stage2_regs_15_0_4 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  stage2_regs_15_0_5 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  stage2_regs_15_0_6 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  stage2_regs_15_0_7 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  stage2_regs_15_0_8 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  stage2_regs_15_1_0 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  stage2_regs_15_1_1 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  stage2_regs_15_1_2 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  stage2_regs_15_1_3 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  stage2_regs_15_1_4 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  stage2_regs_15_1_5 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  stage2_regs_15_1_6 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  stage2_regs_15_1_7 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  stage2_regs_15_1_8 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  stage3_regs_0_0_0 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  stage3_regs_0_0_1 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  stage3_regs_0_0_2 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  stage3_regs_0_0_3 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  stage3_regs_0_0_4 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  stage3_regs_0_0_5 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  stage3_regs_0_0_6 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  stage3_regs_0_0_7 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  stage3_regs_0_0_8 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  stage3_regs_0_0_9 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  stage3_regs_0_0_10 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  stage3_regs_0_0_11 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  stage3_regs_0_1_0 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  stage3_regs_0_1_1 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  stage3_regs_0_1_2 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  stage3_regs_0_1_3 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  stage3_regs_0_1_4 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  stage3_regs_0_1_5 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  stage3_regs_0_1_6 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  stage3_regs_0_1_7 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  stage3_regs_0_1_8 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  stage3_regs_0_1_9 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  stage3_regs_0_1_10 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  stage3_regs_0_1_11 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  stage3_regs_1_0_0 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  stage3_regs_1_0_1 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  stage3_regs_1_0_2 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  stage3_regs_1_0_3 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  stage3_regs_1_0_4 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  stage3_regs_1_0_5 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  stage3_regs_1_0_6 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  stage3_regs_1_0_7 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  stage3_regs_1_0_8 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  stage3_regs_1_0_9 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  stage3_regs_1_0_10 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  stage3_regs_1_0_11 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  stage3_regs_1_1_0 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  stage3_regs_1_1_1 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  stage3_regs_1_1_2 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  stage3_regs_1_1_3 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  stage3_regs_1_1_4 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  stage3_regs_1_1_5 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  stage3_regs_1_1_6 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  stage3_regs_1_1_7 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  stage3_regs_1_1_8 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  stage3_regs_1_1_9 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  stage3_regs_1_1_10 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  stage3_regs_1_1_11 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  stage3_regs_2_0_0 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  stage3_regs_2_0_1 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  stage3_regs_2_0_2 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  stage3_regs_2_0_3 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  stage3_regs_2_0_4 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  stage3_regs_2_0_5 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  stage3_regs_2_0_6 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  stage3_regs_2_0_7 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  stage3_regs_2_0_8 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  stage3_regs_2_0_9 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  stage3_regs_2_0_10 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  stage3_regs_2_0_11 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  stage3_regs_2_1_0 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  stage3_regs_2_1_1 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  stage3_regs_2_1_2 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  stage3_regs_2_1_3 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  stage3_regs_2_1_4 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  stage3_regs_2_1_5 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  stage3_regs_2_1_6 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  stage3_regs_2_1_7 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  stage3_regs_2_1_8 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  stage3_regs_2_1_9 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  stage3_regs_2_1_10 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  stage3_regs_2_1_11 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  stage3_regs_3_0_0 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  stage3_regs_3_0_1 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  stage3_regs_3_0_2 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  stage3_regs_3_0_3 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  stage3_regs_3_0_4 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  stage3_regs_3_0_5 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  stage3_regs_3_0_6 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  stage3_regs_3_0_7 = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  stage3_regs_3_0_8 = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  stage3_regs_3_0_9 = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  stage3_regs_3_0_10 = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  stage3_regs_3_0_11 = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  stage3_regs_3_1_0 = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  stage3_regs_3_1_1 = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  stage3_regs_3_1_2 = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  stage3_regs_3_1_3 = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  stage3_regs_3_1_4 = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  stage3_regs_3_1_5 = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  stage3_regs_3_1_6 = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  stage3_regs_3_1_7 = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  stage3_regs_3_1_8 = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  stage3_regs_3_1_9 = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  stage3_regs_3_1_10 = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  stage3_regs_3_1_11 = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  stage3_regs_4_0_0 = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  stage3_regs_4_0_1 = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  stage3_regs_4_0_2 = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  stage3_regs_4_0_3 = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  stage3_regs_4_0_4 = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  stage3_regs_4_0_5 = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  stage3_regs_4_0_6 = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  stage3_regs_4_0_7 = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  stage3_regs_4_0_8 = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  stage3_regs_4_0_9 = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  stage3_regs_4_0_10 = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  stage3_regs_4_0_11 = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  stage3_regs_4_1_0 = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  stage3_regs_4_1_1 = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  stage3_regs_4_1_2 = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  stage3_regs_4_1_3 = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  stage3_regs_4_1_4 = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  stage3_regs_4_1_5 = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  stage3_regs_4_1_6 = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  stage3_regs_4_1_7 = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  stage3_regs_4_1_8 = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  stage3_regs_4_1_9 = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  stage3_regs_4_1_10 = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  stage3_regs_4_1_11 = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  stage3_regs_5_0_0 = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  stage3_regs_5_0_1 = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  stage3_regs_5_0_2 = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  stage3_regs_5_0_3 = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  stage3_regs_5_0_4 = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  stage3_regs_5_0_5 = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  stage3_regs_5_0_6 = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  stage3_regs_5_0_7 = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  stage3_regs_5_0_8 = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  stage3_regs_5_0_9 = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  stage3_regs_5_0_10 = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  stage3_regs_5_0_11 = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  stage3_regs_5_1_0 = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  stage3_regs_5_1_1 = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  stage3_regs_5_1_2 = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  stage3_regs_5_1_3 = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  stage3_regs_5_1_4 = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  stage3_regs_5_1_5 = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  stage3_regs_5_1_6 = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  stage3_regs_5_1_7 = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  stage3_regs_5_1_8 = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  stage3_regs_5_1_9 = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  stage3_regs_5_1_10 = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  stage3_regs_5_1_11 = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  stage3_regs_6_0_0 = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  stage3_regs_6_0_1 = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  stage3_regs_6_0_2 = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  stage3_regs_6_0_3 = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  stage3_regs_6_0_4 = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  stage3_regs_6_0_5 = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  stage3_regs_6_0_6 = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  stage3_regs_6_0_7 = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  stage3_regs_6_0_8 = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  stage3_regs_6_0_9 = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  stage3_regs_6_0_10 = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  stage3_regs_6_0_11 = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  stage3_regs_6_1_0 = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  stage3_regs_6_1_1 = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  stage3_regs_6_1_2 = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  stage3_regs_6_1_3 = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  stage3_regs_6_1_4 = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  stage3_regs_6_1_5 = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  stage3_regs_6_1_6 = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  stage3_regs_6_1_7 = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  stage3_regs_6_1_8 = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  stage3_regs_6_1_9 = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  stage3_regs_6_1_10 = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  stage3_regs_6_1_11 = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  stage3_regs_7_0_0 = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  stage3_regs_7_0_1 = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  stage3_regs_7_0_2 = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  stage3_regs_7_0_3 = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  stage3_regs_7_0_4 = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  stage3_regs_7_0_5 = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  stage3_regs_7_0_6 = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  stage3_regs_7_0_7 = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  stage3_regs_7_0_8 = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  stage3_regs_7_0_9 = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  stage3_regs_7_0_10 = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  stage3_regs_7_0_11 = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  stage3_regs_7_1_0 = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  stage3_regs_7_1_1 = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  stage3_regs_7_1_2 = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  stage3_regs_7_1_3 = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  stage3_regs_7_1_4 = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  stage3_regs_7_1_5 = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  stage3_regs_7_1_6 = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  stage3_regs_7_1_7 = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  stage3_regs_7_1_8 = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  stage3_regs_7_1_9 = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  stage3_regs_7_1_10 = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  stage3_regs_7_1_11 = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  stage3_regs_8_0_0 = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  stage3_regs_8_0_1 = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  stage3_regs_8_0_2 = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  stage3_regs_8_0_3 = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  stage3_regs_8_0_4 = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  stage3_regs_8_0_5 = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  stage3_regs_8_0_6 = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  stage3_regs_8_0_7 = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  stage3_regs_8_0_8 = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  stage3_regs_8_0_9 = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  stage3_regs_8_0_10 = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  stage3_regs_8_0_11 = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  stage3_regs_8_1_0 = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  stage3_regs_8_1_1 = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  stage3_regs_8_1_2 = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  stage3_regs_8_1_3 = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  stage3_regs_8_1_4 = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  stage3_regs_8_1_5 = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  stage3_regs_8_1_6 = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  stage3_regs_8_1_7 = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  stage3_regs_8_1_8 = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  stage3_regs_8_1_9 = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  stage3_regs_8_1_10 = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  stage3_regs_8_1_11 = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  stage3_regs_9_0_0 = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  stage3_regs_9_0_1 = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  stage3_regs_9_0_2 = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  stage3_regs_9_0_3 = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  stage3_regs_9_0_4 = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  stage3_regs_9_0_5 = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  stage3_regs_9_0_6 = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  stage3_regs_9_0_7 = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  stage3_regs_9_0_8 = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  stage3_regs_9_0_9 = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  stage3_regs_9_0_10 = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  stage3_regs_9_0_11 = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  stage3_regs_9_1_0 = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  stage3_regs_9_1_1 = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  stage3_regs_9_1_2 = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  stage3_regs_9_1_3 = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  stage3_regs_9_1_4 = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  stage3_regs_9_1_5 = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  stage3_regs_9_1_6 = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  stage3_regs_9_1_7 = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  stage3_regs_9_1_8 = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  stage3_regs_9_1_9 = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  stage3_regs_9_1_10 = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  stage3_regs_9_1_11 = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  stage3_regs_10_0_0 = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  stage3_regs_10_0_1 = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  stage3_regs_10_0_2 = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  stage3_regs_10_0_3 = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  stage3_regs_10_0_4 = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  stage3_regs_10_0_5 = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  stage3_regs_10_0_6 = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  stage3_regs_10_0_7 = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  stage3_regs_10_0_8 = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  stage3_regs_10_0_9 = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  stage3_regs_10_0_10 = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  stage3_regs_10_0_11 = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  stage3_regs_10_1_0 = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  stage3_regs_10_1_1 = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  stage3_regs_10_1_2 = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  stage3_regs_10_1_3 = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  stage3_regs_10_1_4 = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  stage3_regs_10_1_5 = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  stage3_regs_10_1_6 = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  stage3_regs_10_1_7 = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  stage3_regs_10_1_8 = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  stage3_regs_10_1_9 = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  stage3_regs_10_1_10 = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  stage3_regs_10_1_11 = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  stage3_regs_11_0_0 = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  stage3_regs_11_0_1 = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  stage3_regs_11_0_2 = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  stage3_regs_11_0_3 = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  stage3_regs_11_0_4 = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  stage3_regs_11_0_5 = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  stage3_regs_11_0_6 = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  stage3_regs_11_0_7 = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  stage3_regs_11_0_8 = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  stage3_regs_11_0_9 = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  stage3_regs_11_0_10 = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  stage3_regs_11_0_11 = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  stage3_regs_11_1_0 = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  stage3_regs_11_1_1 = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  stage3_regs_11_1_2 = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  stage3_regs_11_1_3 = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  stage3_regs_11_1_4 = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  stage3_regs_11_1_5 = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  stage3_regs_11_1_6 = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  stage3_regs_11_1_7 = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  stage3_regs_11_1_8 = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  stage3_regs_11_1_9 = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  stage3_regs_11_1_10 = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  stage3_regs_11_1_11 = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  stage3_regs_12_0_0 = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  stage3_regs_12_0_1 = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  stage3_regs_12_0_2 = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  stage3_regs_12_0_3 = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  stage3_regs_12_0_4 = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  stage3_regs_12_0_5 = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  stage3_regs_12_0_6 = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  stage3_regs_12_0_7 = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  stage3_regs_12_0_8 = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  stage3_regs_12_0_9 = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  stage3_regs_12_0_10 = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  stage3_regs_12_0_11 = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  stage3_regs_12_1_0 = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  stage3_regs_12_1_1 = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  stage3_regs_12_1_2 = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  stage3_regs_12_1_3 = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  stage3_regs_12_1_4 = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  stage3_regs_12_1_5 = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  stage3_regs_12_1_6 = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  stage3_regs_12_1_7 = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  stage3_regs_12_1_8 = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  stage3_regs_12_1_9 = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  stage3_regs_12_1_10 = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  stage3_regs_12_1_11 = _RAND_999[31:0];
  _RAND_1000 = {1{`RANDOM}};
  stage3_regs_13_0_0 = _RAND_1000[31:0];
  _RAND_1001 = {1{`RANDOM}};
  stage3_regs_13_0_1 = _RAND_1001[31:0];
  _RAND_1002 = {1{`RANDOM}};
  stage3_regs_13_0_2 = _RAND_1002[31:0];
  _RAND_1003 = {1{`RANDOM}};
  stage3_regs_13_0_3 = _RAND_1003[31:0];
  _RAND_1004 = {1{`RANDOM}};
  stage3_regs_13_0_4 = _RAND_1004[31:0];
  _RAND_1005 = {1{`RANDOM}};
  stage3_regs_13_0_5 = _RAND_1005[31:0];
  _RAND_1006 = {1{`RANDOM}};
  stage3_regs_13_0_6 = _RAND_1006[31:0];
  _RAND_1007 = {1{`RANDOM}};
  stage3_regs_13_0_7 = _RAND_1007[31:0];
  _RAND_1008 = {1{`RANDOM}};
  stage3_regs_13_0_8 = _RAND_1008[31:0];
  _RAND_1009 = {1{`RANDOM}};
  stage3_regs_13_0_9 = _RAND_1009[31:0];
  _RAND_1010 = {1{`RANDOM}};
  stage3_regs_13_0_10 = _RAND_1010[31:0];
  _RAND_1011 = {1{`RANDOM}};
  stage3_regs_13_0_11 = _RAND_1011[31:0];
  _RAND_1012 = {1{`RANDOM}};
  stage3_regs_13_1_0 = _RAND_1012[31:0];
  _RAND_1013 = {1{`RANDOM}};
  stage3_regs_13_1_1 = _RAND_1013[31:0];
  _RAND_1014 = {1{`RANDOM}};
  stage3_regs_13_1_2 = _RAND_1014[31:0];
  _RAND_1015 = {1{`RANDOM}};
  stage3_regs_13_1_3 = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  stage3_regs_13_1_4 = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  stage3_regs_13_1_5 = _RAND_1017[31:0];
  _RAND_1018 = {1{`RANDOM}};
  stage3_regs_13_1_6 = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  stage3_regs_13_1_7 = _RAND_1019[31:0];
  _RAND_1020 = {1{`RANDOM}};
  stage3_regs_13_1_8 = _RAND_1020[31:0];
  _RAND_1021 = {1{`RANDOM}};
  stage3_regs_13_1_9 = _RAND_1021[31:0];
  _RAND_1022 = {1{`RANDOM}};
  stage3_regs_13_1_10 = _RAND_1022[31:0];
  _RAND_1023 = {1{`RANDOM}};
  stage3_regs_13_1_11 = _RAND_1023[31:0];
  _RAND_1024 = {1{`RANDOM}};
  stage3_regs_14_0_0 = _RAND_1024[31:0];
  _RAND_1025 = {1{`RANDOM}};
  stage3_regs_14_0_1 = _RAND_1025[31:0];
  _RAND_1026 = {1{`RANDOM}};
  stage3_regs_14_0_2 = _RAND_1026[31:0];
  _RAND_1027 = {1{`RANDOM}};
  stage3_regs_14_0_3 = _RAND_1027[31:0];
  _RAND_1028 = {1{`RANDOM}};
  stage3_regs_14_0_4 = _RAND_1028[31:0];
  _RAND_1029 = {1{`RANDOM}};
  stage3_regs_14_0_5 = _RAND_1029[31:0];
  _RAND_1030 = {1{`RANDOM}};
  stage3_regs_14_0_6 = _RAND_1030[31:0];
  _RAND_1031 = {1{`RANDOM}};
  stage3_regs_14_0_7 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  stage3_regs_14_0_8 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  stage3_regs_14_0_9 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  stage3_regs_14_0_10 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  stage3_regs_14_0_11 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  stage3_regs_14_1_0 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  stage3_regs_14_1_1 = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  stage3_regs_14_1_2 = _RAND_1038[31:0];
  _RAND_1039 = {1{`RANDOM}};
  stage3_regs_14_1_3 = _RAND_1039[31:0];
  _RAND_1040 = {1{`RANDOM}};
  stage3_regs_14_1_4 = _RAND_1040[31:0];
  _RAND_1041 = {1{`RANDOM}};
  stage3_regs_14_1_5 = _RAND_1041[31:0];
  _RAND_1042 = {1{`RANDOM}};
  stage3_regs_14_1_6 = _RAND_1042[31:0];
  _RAND_1043 = {1{`RANDOM}};
  stage3_regs_14_1_7 = _RAND_1043[31:0];
  _RAND_1044 = {1{`RANDOM}};
  stage3_regs_14_1_8 = _RAND_1044[31:0];
  _RAND_1045 = {1{`RANDOM}};
  stage3_regs_14_1_9 = _RAND_1045[31:0];
  _RAND_1046 = {1{`RANDOM}};
  stage3_regs_14_1_10 = _RAND_1046[31:0];
  _RAND_1047 = {1{`RANDOM}};
  stage3_regs_14_1_11 = _RAND_1047[31:0];
  _RAND_1048 = {1{`RANDOM}};
  stage3_regs_15_0_0 = _RAND_1048[31:0];
  _RAND_1049 = {1{`RANDOM}};
  stage3_regs_15_0_1 = _RAND_1049[31:0];
  _RAND_1050 = {1{`RANDOM}};
  stage3_regs_15_0_2 = _RAND_1050[31:0];
  _RAND_1051 = {1{`RANDOM}};
  stage3_regs_15_0_3 = _RAND_1051[31:0];
  _RAND_1052 = {1{`RANDOM}};
  stage3_regs_15_0_4 = _RAND_1052[31:0];
  _RAND_1053 = {1{`RANDOM}};
  stage3_regs_15_0_5 = _RAND_1053[31:0];
  _RAND_1054 = {1{`RANDOM}};
  stage3_regs_15_0_6 = _RAND_1054[31:0];
  _RAND_1055 = {1{`RANDOM}};
  stage3_regs_15_0_7 = _RAND_1055[31:0];
  _RAND_1056 = {1{`RANDOM}};
  stage3_regs_15_0_8 = _RAND_1056[31:0];
  _RAND_1057 = {1{`RANDOM}};
  stage3_regs_15_0_9 = _RAND_1057[31:0];
  _RAND_1058 = {1{`RANDOM}};
  stage3_regs_15_0_10 = _RAND_1058[31:0];
  _RAND_1059 = {1{`RANDOM}};
  stage3_regs_15_0_11 = _RAND_1059[31:0];
  _RAND_1060 = {1{`RANDOM}};
  stage3_regs_15_1_0 = _RAND_1060[31:0];
  _RAND_1061 = {1{`RANDOM}};
  stage3_regs_15_1_1 = _RAND_1061[31:0];
  _RAND_1062 = {1{`RANDOM}};
  stage3_regs_15_1_2 = _RAND_1062[31:0];
  _RAND_1063 = {1{`RANDOM}};
  stage3_regs_15_1_3 = _RAND_1063[31:0];
  _RAND_1064 = {1{`RANDOM}};
  stage3_regs_15_1_4 = _RAND_1064[31:0];
  _RAND_1065 = {1{`RANDOM}};
  stage3_regs_15_1_5 = _RAND_1065[31:0];
  _RAND_1066 = {1{`RANDOM}};
  stage3_regs_15_1_6 = _RAND_1066[31:0];
  _RAND_1067 = {1{`RANDOM}};
  stage3_regs_15_1_7 = _RAND_1067[31:0];
  _RAND_1068 = {1{`RANDOM}};
  stage3_regs_15_1_8 = _RAND_1068[31:0];
  _RAND_1069 = {1{`RANDOM}};
  stage3_regs_15_1_9 = _RAND_1069[31:0];
  _RAND_1070 = {1{`RANDOM}};
  stage3_regs_15_1_10 = _RAND_1070[31:0];
  _RAND_1071 = {1{`RANDOM}};
  stage3_regs_15_1_11 = _RAND_1071[31:0];
  _RAND_1072 = {1{`RANDOM}};
  stage4_regs_0_1_0 = _RAND_1072[31:0];
  _RAND_1073 = {1{`RANDOM}};
  stage4_regs_0_1_1 = _RAND_1073[31:0];
  _RAND_1074 = {1{`RANDOM}};
  stage4_regs_0_1_2 = _RAND_1074[31:0];
  _RAND_1075 = {1{`RANDOM}};
  stage4_regs_0_1_3 = _RAND_1075[31:0];
  _RAND_1076 = {1{`RANDOM}};
  stage4_regs_0_1_4 = _RAND_1076[31:0];
  _RAND_1077 = {1{`RANDOM}};
  stage4_regs_0_1_5 = _RAND_1077[31:0];
  _RAND_1078 = {1{`RANDOM}};
  stage4_regs_0_1_6 = _RAND_1078[31:0];
  _RAND_1079 = {1{`RANDOM}};
  stage4_regs_0_1_7 = _RAND_1079[31:0];
  _RAND_1080 = {1{`RANDOM}};
  stage4_regs_0_1_8 = _RAND_1080[31:0];
  _RAND_1081 = {1{`RANDOM}};
  stage4_regs_1_1_0 = _RAND_1081[31:0];
  _RAND_1082 = {1{`RANDOM}};
  stage4_regs_1_1_1 = _RAND_1082[31:0];
  _RAND_1083 = {1{`RANDOM}};
  stage4_regs_1_1_2 = _RAND_1083[31:0];
  _RAND_1084 = {1{`RANDOM}};
  stage4_regs_1_1_3 = _RAND_1084[31:0];
  _RAND_1085 = {1{`RANDOM}};
  stage4_regs_1_1_4 = _RAND_1085[31:0];
  _RAND_1086 = {1{`RANDOM}};
  stage4_regs_1_1_5 = _RAND_1086[31:0];
  _RAND_1087 = {1{`RANDOM}};
  stage4_regs_1_1_6 = _RAND_1087[31:0];
  _RAND_1088 = {1{`RANDOM}};
  stage4_regs_1_1_7 = _RAND_1088[31:0];
  _RAND_1089 = {1{`RANDOM}};
  stage4_regs_1_1_8 = _RAND_1089[31:0];
  _RAND_1090 = {1{`RANDOM}};
  stage4_regs_2_1_0 = _RAND_1090[31:0];
  _RAND_1091 = {1{`RANDOM}};
  stage4_regs_2_1_1 = _RAND_1091[31:0];
  _RAND_1092 = {1{`RANDOM}};
  stage4_regs_2_1_2 = _RAND_1092[31:0];
  _RAND_1093 = {1{`RANDOM}};
  stage4_regs_2_1_3 = _RAND_1093[31:0];
  _RAND_1094 = {1{`RANDOM}};
  stage4_regs_2_1_4 = _RAND_1094[31:0];
  _RAND_1095 = {1{`RANDOM}};
  stage4_regs_2_1_5 = _RAND_1095[31:0];
  _RAND_1096 = {1{`RANDOM}};
  stage4_regs_2_1_6 = _RAND_1096[31:0];
  _RAND_1097 = {1{`RANDOM}};
  stage4_regs_2_1_7 = _RAND_1097[31:0];
  _RAND_1098 = {1{`RANDOM}};
  stage4_regs_2_1_8 = _RAND_1098[31:0];
  _RAND_1099 = {1{`RANDOM}};
  stage4_regs_3_1_0 = _RAND_1099[31:0];
  _RAND_1100 = {1{`RANDOM}};
  stage4_regs_3_1_1 = _RAND_1100[31:0];
  _RAND_1101 = {1{`RANDOM}};
  stage4_regs_3_1_2 = _RAND_1101[31:0];
  _RAND_1102 = {1{`RANDOM}};
  stage4_regs_3_1_3 = _RAND_1102[31:0];
  _RAND_1103 = {1{`RANDOM}};
  stage4_regs_3_1_4 = _RAND_1103[31:0];
  _RAND_1104 = {1{`RANDOM}};
  stage4_regs_3_1_5 = _RAND_1104[31:0];
  _RAND_1105 = {1{`RANDOM}};
  stage4_regs_3_1_6 = _RAND_1105[31:0];
  _RAND_1106 = {1{`RANDOM}};
  stage4_regs_3_1_7 = _RAND_1106[31:0];
  _RAND_1107 = {1{`RANDOM}};
  stage4_regs_3_1_8 = _RAND_1107[31:0];
  _RAND_1108 = {1{`RANDOM}};
  stage4_regs_4_1_0 = _RAND_1108[31:0];
  _RAND_1109 = {1{`RANDOM}};
  stage4_regs_4_1_1 = _RAND_1109[31:0];
  _RAND_1110 = {1{`RANDOM}};
  stage4_regs_4_1_2 = _RAND_1110[31:0];
  _RAND_1111 = {1{`RANDOM}};
  stage4_regs_4_1_3 = _RAND_1111[31:0];
  _RAND_1112 = {1{`RANDOM}};
  stage4_regs_4_1_4 = _RAND_1112[31:0];
  _RAND_1113 = {1{`RANDOM}};
  stage4_regs_4_1_5 = _RAND_1113[31:0];
  _RAND_1114 = {1{`RANDOM}};
  stage4_regs_4_1_6 = _RAND_1114[31:0];
  _RAND_1115 = {1{`RANDOM}};
  stage4_regs_4_1_7 = _RAND_1115[31:0];
  _RAND_1116 = {1{`RANDOM}};
  stage4_regs_4_1_8 = _RAND_1116[31:0];
  _RAND_1117 = {1{`RANDOM}};
  stage4_regs_5_1_0 = _RAND_1117[31:0];
  _RAND_1118 = {1{`RANDOM}};
  stage4_regs_5_1_1 = _RAND_1118[31:0];
  _RAND_1119 = {1{`RANDOM}};
  stage4_regs_5_1_2 = _RAND_1119[31:0];
  _RAND_1120 = {1{`RANDOM}};
  stage4_regs_5_1_3 = _RAND_1120[31:0];
  _RAND_1121 = {1{`RANDOM}};
  stage4_regs_5_1_4 = _RAND_1121[31:0];
  _RAND_1122 = {1{`RANDOM}};
  stage4_regs_5_1_5 = _RAND_1122[31:0];
  _RAND_1123 = {1{`RANDOM}};
  stage4_regs_5_1_6 = _RAND_1123[31:0];
  _RAND_1124 = {1{`RANDOM}};
  stage4_regs_5_1_7 = _RAND_1124[31:0];
  _RAND_1125 = {1{`RANDOM}};
  stage4_regs_5_1_8 = _RAND_1125[31:0];
  _RAND_1126 = {1{`RANDOM}};
  stage4_regs_6_1_0 = _RAND_1126[31:0];
  _RAND_1127 = {1{`RANDOM}};
  stage4_regs_6_1_1 = _RAND_1127[31:0];
  _RAND_1128 = {1{`RANDOM}};
  stage4_regs_6_1_2 = _RAND_1128[31:0];
  _RAND_1129 = {1{`RANDOM}};
  stage4_regs_6_1_3 = _RAND_1129[31:0];
  _RAND_1130 = {1{`RANDOM}};
  stage4_regs_6_1_4 = _RAND_1130[31:0];
  _RAND_1131 = {1{`RANDOM}};
  stage4_regs_6_1_5 = _RAND_1131[31:0];
  _RAND_1132 = {1{`RANDOM}};
  stage4_regs_6_1_6 = _RAND_1132[31:0];
  _RAND_1133 = {1{`RANDOM}};
  stage4_regs_6_1_7 = _RAND_1133[31:0];
  _RAND_1134 = {1{`RANDOM}};
  stage4_regs_6_1_8 = _RAND_1134[31:0];
  _RAND_1135 = {1{`RANDOM}};
  stage4_regs_7_1_0 = _RAND_1135[31:0];
  _RAND_1136 = {1{`RANDOM}};
  stage4_regs_7_1_1 = _RAND_1136[31:0];
  _RAND_1137 = {1{`RANDOM}};
  stage4_regs_7_1_2 = _RAND_1137[31:0];
  _RAND_1138 = {1{`RANDOM}};
  stage4_regs_7_1_3 = _RAND_1138[31:0];
  _RAND_1139 = {1{`RANDOM}};
  stage4_regs_7_1_4 = _RAND_1139[31:0];
  _RAND_1140 = {1{`RANDOM}};
  stage4_regs_7_1_5 = _RAND_1140[31:0];
  _RAND_1141 = {1{`RANDOM}};
  stage4_regs_7_1_6 = _RAND_1141[31:0];
  _RAND_1142 = {1{`RANDOM}};
  stage4_regs_7_1_7 = _RAND_1142[31:0];
  _RAND_1143 = {1{`RANDOM}};
  stage4_regs_7_1_8 = _RAND_1143[31:0];
  _RAND_1144 = {1{`RANDOM}};
  stage4_regs_8_1_0 = _RAND_1144[31:0];
  _RAND_1145 = {1{`RANDOM}};
  stage4_regs_8_1_1 = _RAND_1145[31:0];
  _RAND_1146 = {1{`RANDOM}};
  stage4_regs_8_1_2 = _RAND_1146[31:0];
  _RAND_1147 = {1{`RANDOM}};
  stage4_regs_8_1_3 = _RAND_1147[31:0];
  _RAND_1148 = {1{`RANDOM}};
  stage4_regs_8_1_4 = _RAND_1148[31:0];
  _RAND_1149 = {1{`RANDOM}};
  stage4_regs_8_1_5 = _RAND_1149[31:0];
  _RAND_1150 = {1{`RANDOM}};
  stage4_regs_8_1_6 = _RAND_1150[31:0];
  _RAND_1151 = {1{`RANDOM}};
  stage4_regs_8_1_7 = _RAND_1151[31:0];
  _RAND_1152 = {1{`RANDOM}};
  stage4_regs_8_1_8 = _RAND_1152[31:0];
  _RAND_1153 = {1{`RANDOM}};
  stage4_regs_9_1_0 = _RAND_1153[31:0];
  _RAND_1154 = {1{`RANDOM}};
  stage4_regs_9_1_1 = _RAND_1154[31:0];
  _RAND_1155 = {1{`RANDOM}};
  stage4_regs_9_1_2 = _RAND_1155[31:0];
  _RAND_1156 = {1{`RANDOM}};
  stage4_regs_9_1_3 = _RAND_1156[31:0];
  _RAND_1157 = {1{`RANDOM}};
  stage4_regs_9_1_4 = _RAND_1157[31:0];
  _RAND_1158 = {1{`RANDOM}};
  stage4_regs_9_1_5 = _RAND_1158[31:0];
  _RAND_1159 = {1{`RANDOM}};
  stage4_regs_9_1_6 = _RAND_1159[31:0];
  _RAND_1160 = {1{`RANDOM}};
  stage4_regs_9_1_7 = _RAND_1160[31:0];
  _RAND_1161 = {1{`RANDOM}};
  stage4_regs_9_1_8 = _RAND_1161[31:0];
  _RAND_1162 = {1{`RANDOM}};
  stage4_regs_10_1_0 = _RAND_1162[31:0];
  _RAND_1163 = {1{`RANDOM}};
  stage4_regs_10_1_1 = _RAND_1163[31:0];
  _RAND_1164 = {1{`RANDOM}};
  stage4_regs_10_1_2 = _RAND_1164[31:0];
  _RAND_1165 = {1{`RANDOM}};
  stage4_regs_10_1_3 = _RAND_1165[31:0];
  _RAND_1166 = {1{`RANDOM}};
  stage4_regs_10_1_4 = _RAND_1166[31:0];
  _RAND_1167 = {1{`RANDOM}};
  stage4_regs_10_1_5 = _RAND_1167[31:0];
  _RAND_1168 = {1{`RANDOM}};
  stage4_regs_10_1_6 = _RAND_1168[31:0];
  _RAND_1169 = {1{`RANDOM}};
  stage4_regs_10_1_7 = _RAND_1169[31:0];
  _RAND_1170 = {1{`RANDOM}};
  stage4_regs_10_1_8 = _RAND_1170[31:0];
  _RAND_1171 = {1{`RANDOM}};
  stage4_regs_11_1_0 = _RAND_1171[31:0];
  _RAND_1172 = {1{`RANDOM}};
  stage4_regs_11_1_1 = _RAND_1172[31:0];
  _RAND_1173 = {1{`RANDOM}};
  stage4_regs_11_1_2 = _RAND_1173[31:0];
  _RAND_1174 = {1{`RANDOM}};
  stage4_regs_11_1_3 = _RAND_1174[31:0];
  _RAND_1175 = {1{`RANDOM}};
  stage4_regs_11_1_4 = _RAND_1175[31:0];
  _RAND_1176 = {1{`RANDOM}};
  stage4_regs_11_1_5 = _RAND_1176[31:0];
  _RAND_1177 = {1{`RANDOM}};
  stage4_regs_11_1_6 = _RAND_1177[31:0];
  _RAND_1178 = {1{`RANDOM}};
  stage4_regs_11_1_7 = _RAND_1178[31:0];
  _RAND_1179 = {1{`RANDOM}};
  stage4_regs_11_1_8 = _RAND_1179[31:0];
  _RAND_1180 = {1{`RANDOM}};
  stage4_regs_12_1_0 = _RAND_1180[31:0];
  _RAND_1181 = {1{`RANDOM}};
  stage4_regs_12_1_1 = _RAND_1181[31:0];
  _RAND_1182 = {1{`RANDOM}};
  stage4_regs_12_1_2 = _RAND_1182[31:0];
  _RAND_1183 = {1{`RANDOM}};
  stage4_regs_12_1_3 = _RAND_1183[31:0];
  _RAND_1184 = {1{`RANDOM}};
  stage4_regs_12_1_4 = _RAND_1184[31:0];
  _RAND_1185 = {1{`RANDOM}};
  stage4_regs_12_1_5 = _RAND_1185[31:0];
  _RAND_1186 = {1{`RANDOM}};
  stage4_regs_12_1_6 = _RAND_1186[31:0];
  _RAND_1187 = {1{`RANDOM}};
  stage4_regs_12_1_7 = _RAND_1187[31:0];
  _RAND_1188 = {1{`RANDOM}};
  stage4_regs_12_1_8 = _RAND_1188[31:0];
  _RAND_1189 = {1{`RANDOM}};
  stage4_regs_13_1_0 = _RAND_1189[31:0];
  _RAND_1190 = {1{`RANDOM}};
  stage4_regs_13_1_1 = _RAND_1190[31:0];
  _RAND_1191 = {1{`RANDOM}};
  stage4_regs_13_1_2 = _RAND_1191[31:0];
  _RAND_1192 = {1{`RANDOM}};
  stage4_regs_13_1_3 = _RAND_1192[31:0];
  _RAND_1193 = {1{`RANDOM}};
  stage4_regs_13_1_4 = _RAND_1193[31:0];
  _RAND_1194 = {1{`RANDOM}};
  stage4_regs_13_1_5 = _RAND_1194[31:0];
  _RAND_1195 = {1{`RANDOM}};
  stage4_regs_13_1_6 = _RAND_1195[31:0];
  _RAND_1196 = {1{`RANDOM}};
  stage4_regs_13_1_7 = _RAND_1196[31:0];
  _RAND_1197 = {1{`RANDOM}};
  stage4_regs_13_1_8 = _RAND_1197[31:0];
  _RAND_1198 = {1{`RANDOM}};
  stage4_regs_14_1_0 = _RAND_1198[31:0];
  _RAND_1199 = {1{`RANDOM}};
  stage4_regs_14_1_1 = _RAND_1199[31:0];
  _RAND_1200 = {1{`RANDOM}};
  stage4_regs_14_1_2 = _RAND_1200[31:0];
  _RAND_1201 = {1{`RANDOM}};
  stage4_regs_14_1_3 = _RAND_1201[31:0];
  _RAND_1202 = {1{`RANDOM}};
  stage4_regs_14_1_4 = _RAND_1202[31:0];
  _RAND_1203 = {1{`RANDOM}};
  stage4_regs_14_1_5 = _RAND_1203[31:0];
  _RAND_1204 = {1{`RANDOM}};
  stage4_regs_14_1_6 = _RAND_1204[31:0];
  _RAND_1205 = {1{`RANDOM}};
  stage4_regs_14_1_7 = _RAND_1205[31:0];
  _RAND_1206 = {1{`RANDOM}};
  stage4_regs_14_1_8 = _RAND_1206[31:0];
  _RAND_1207 = {1{`RANDOM}};
  stage4_regs_15_1_0 = _RAND_1207[31:0];
  _RAND_1208 = {1{`RANDOM}};
  stage4_regs_15_1_1 = _RAND_1208[31:0];
  _RAND_1209 = {1{`RANDOM}};
  stage4_regs_15_1_2 = _RAND_1209[31:0];
  _RAND_1210 = {1{`RANDOM}};
  stage4_regs_15_1_3 = _RAND_1210[31:0];
  _RAND_1211 = {1{`RANDOM}};
  stage4_regs_15_1_4 = _RAND_1211[31:0];
  _RAND_1212 = {1{`RANDOM}};
  stage4_regs_15_1_5 = _RAND_1212[31:0];
  _RAND_1213 = {1{`RANDOM}};
  stage4_regs_15_1_6 = _RAND_1213[31:0];
  _RAND_1214 = {1{`RANDOM}};
  stage4_regs_15_1_7 = _RAND_1214[31:0];
  _RAND_1215 = {1{`RANDOM}};
  stage4_regs_15_1_8 = _RAND_1215[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPU_hs_lib(
  input         clock,
  input         reset,
  input         io_add_en,
  input  [31:0] io_add_a,
  input  [31:0] io_add_b,
  output [31:0] io_add_s,
  input         io_sub_en,
  input  [31:0] io_sub_a,
  input  [31:0] io_sub_b,
  output [31:0] io_sub_s,
  input         io_mul_en,
  input  [31:0] io_mul_a,
  input  [31:0] io_mul_b,
  output [31:0] io_mul_s,
  input         io_div_en,
  input  [31:0] io_div_a,
  input  [31:0] io_div_b,
  output [31:0] io_div_s,
  input         io_rec_en,
  input  [31:0] io_rec_a,
  output [31:0] io_rec_s,
  input         io_sqr_en,
  input  [31:0] io_sqr_a,
  output [31:0] io_sqr_s
);
  wire  FP_adder_13ccs_clock; // @[FloatingPointDesigns.scala 39:21]
  wire  FP_adder_13ccs_reset; // @[FloatingPointDesigns.scala 39:21]
  wire  FP_adder_13ccs_io_in_en; // @[FloatingPointDesigns.scala 39:21]
  wire [31:0] FP_adder_13ccs_io_in_a; // @[FloatingPointDesigns.scala 39:21]
  wire [31:0] FP_adder_13ccs_io_in_b; // @[FloatingPointDesigns.scala 39:21]
  wire [31:0] FP_adder_13ccs_io_out_s; // @[FloatingPointDesigns.scala 39:21]
  wire  FP_subtractor_13ccs_clock; // @[FloatingPointDesigns.scala 40:21]
  wire  FP_subtractor_13ccs_reset; // @[FloatingPointDesigns.scala 40:21]
  wire  FP_subtractor_13ccs_io_in_en; // @[FloatingPointDesigns.scala 40:21]
  wire [31:0] FP_subtractor_13ccs_io_in_a; // @[FloatingPointDesigns.scala 40:21]
  wire [31:0] FP_subtractor_13ccs_io_in_b; // @[FloatingPointDesigns.scala 40:21]
  wire [31:0] FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 40:21]
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 41:21]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 41:21]
  wire  FP_multiplier_10ccs_io_in_en; // @[FloatingPointDesigns.scala 41:21]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 41:21]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 41:21]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 41:21]
  wire  FP_reciprocal_newfpu_clock; // @[FloatingPointDesigns.scala 42:21]
  wire  FP_reciprocal_newfpu_reset; // @[FloatingPointDesigns.scala 42:21]
  wire  FP_reciprocal_newfpu_io_in_en; // @[FloatingPointDesigns.scala 42:21]
  wire [31:0] FP_reciprocal_newfpu_io_in_a; // @[FloatingPointDesigns.scala 42:21]
  wire [31:0] FP_reciprocal_newfpu_io_out_s; // @[FloatingPointDesigns.scala 42:21]
  wire  FP_divider_newfpu_clock; // @[FloatingPointDesigns.scala 43:21]
  wire  FP_divider_newfpu_reset; // @[FloatingPointDesigns.scala 43:21]
  wire  FP_divider_newfpu_io_in_en; // @[FloatingPointDesigns.scala 43:21]
  wire [31:0] FP_divider_newfpu_io_in_a; // @[FloatingPointDesigns.scala 43:21]
  wire [31:0] FP_divider_newfpu_io_in_b; // @[FloatingPointDesigns.scala 43:21]
  wire [31:0] FP_divider_newfpu_io_out_s; // @[FloatingPointDesigns.scala 43:21]
  wire  FP_square_root_newfpu_clock; // @[FloatingPointDesigns.scala 44:21]
  wire  FP_square_root_newfpu_reset; // @[FloatingPointDesigns.scala 44:21]
  wire  FP_square_root_newfpu_io_in_en; // @[FloatingPointDesigns.scala 44:21]
  wire [31:0] FP_square_root_newfpu_io_in_a; // @[FloatingPointDesigns.scala 44:21]
  wire [31:0] FP_square_root_newfpu_io_out_s; // @[FloatingPointDesigns.scala 44:21]
  FP_adder_13ccs FP_adder_13ccs ( // @[FloatingPointDesigns.scala 39:21]
    .clock(FP_adder_13ccs_clock),
    .reset(FP_adder_13ccs_reset),
    .io_in_en(FP_adder_13ccs_io_in_en),
    .io_in_a(FP_adder_13ccs_io_in_a),
    .io_in_b(FP_adder_13ccs_io_in_b),
    .io_out_s(FP_adder_13ccs_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs ( // @[FloatingPointDesigns.scala 40:21]
    .clock(FP_subtractor_13ccs_clock),
    .reset(FP_subtractor_13ccs_reset),
    .io_in_en(FP_subtractor_13ccs_io_in_en),
    .io_in_a(FP_subtractor_13ccs_io_in_a),
    .io_in_b(FP_subtractor_13ccs_io_in_b),
    .io_out_s(FP_subtractor_13ccs_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 41:21]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_en(FP_multiplier_10ccs_io_in_en),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  FP_reciprocal_newfpu FP_reciprocal_newfpu ( // @[FloatingPointDesigns.scala 42:21]
    .clock(FP_reciprocal_newfpu_clock),
    .reset(FP_reciprocal_newfpu_reset),
    .io_in_en(FP_reciprocal_newfpu_io_in_en),
    .io_in_a(FP_reciprocal_newfpu_io_in_a),
    .io_out_s(FP_reciprocal_newfpu_io_out_s)
  );
  FP_divider_newfpu FP_divider_newfpu ( // @[FloatingPointDesigns.scala 43:21]
    .clock(FP_divider_newfpu_clock),
    .reset(FP_divider_newfpu_reset),
    .io_in_en(FP_divider_newfpu_io_in_en),
    .io_in_a(FP_divider_newfpu_io_in_a),
    .io_in_b(FP_divider_newfpu_io_in_b),
    .io_out_s(FP_divider_newfpu_io_out_s)
  );
  FP_square_root_newfpu FP_square_root_newfpu ( // @[FloatingPointDesigns.scala 44:21]
    .clock(FP_square_root_newfpu_clock),
    .reset(FP_square_root_newfpu_reset),
    .io_in_en(FP_square_root_newfpu_io_in_en),
    .io_in_a(FP_square_root_newfpu_io_in_a),
    .io_out_s(FP_square_root_newfpu_io_out_s)
  );
  assign io_add_s = FP_adder_13ccs_io_out_s; // @[FloatingPointDesigns.scala 48:14]
  assign io_sub_s = FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 52:14]
  assign io_mul_s = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 56:14]
  assign io_div_s = FP_divider_newfpu_io_out_s; // @[FloatingPointDesigns.scala 60:14]
  assign io_rec_s = FP_reciprocal_newfpu_io_out_s; // @[FloatingPointDesigns.scala 63:14]
  assign io_sqr_s = FP_square_root_newfpu_io_out_s; // @[FloatingPointDesigns.scala 66:14]
  assign FP_adder_13ccs_clock = clock;
  assign FP_adder_13ccs_reset = reset;
  assign FP_adder_13ccs_io_in_en = io_add_en; // @[FloatingPointDesigns.scala 45:14]
  assign FP_adder_13ccs_io_in_a = io_add_a; // @[FloatingPointDesigns.scala 46:14]
  assign FP_adder_13ccs_io_in_b = io_add_b; // @[FloatingPointDesigns.scala 47:14]
  assign FP_subtractor_13ccs_clock = clock;
  assign FP_subtractor_13ccs_reset = reset;
  assign FP_subtractor_13ccs_io_in_en = io_sub_en; // @[FloatingPointDesigns.scala 49:14]
  assign FP_subtractor_13ccs_io_in_a = io_sub_a; // @[FloatingPointDesigns.scala 50:14]
  assign FP_subtractor_13ccs_io_in_b = io_sub_b; // @[FloatingPointDesigns.scala 51:14]
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_en = io_mul_en; // @[FloatingPointDesigns.scala 53:14]
  assign FP_multiplier_10ccs_io_in_a = io_mul_a; // @[FloatingPointDesigns.scala 54:14]
  assign FP_multiplier_10ccs_io_in_b = io_mul_b; // @[FloatingPointDesigns.scala 55:14]
  assign FP_reciprocal_newfpu_clock = clock;
  assign FP_reciprocal_newfpu_reset = reset;
  assign FP_reciprocal_newfpu_io_in_en = io_rec_en; // @[FloatingPointDesigns.scala 61:14]
  assign FP_reciprocal_newfpu_io_in_a = io_rec_a; // @[FloatingPointDesigns.scala 62:14]
  assign FP_divider_newfpu_clock = clock;
  assign FP_divider_newfpu_reset = reset;
  assign FP_divider_newfpu_io_in_en = io_div_en; // @[FloatingPointDesigns.scala 57:14]
  assign FP_divider_newfpu_io_in_a = io_div_a; // @[FloatingPointDesigns.scala 58:14]
  assign FP_divider_newfpu_io_in_b = io_div_b; // @[FloatingPointDesigns.scala 59:14]
  assign FP_square_root_newfpu_clock = clock;
  assign FP_square_root_newfpu_reset = reset;
  assign FP_square_root_newfpu_io_in_en = io_sqr_en; // @[FloatingPointDesigns.scala 64:14]
  assign FP_square_root_newfpu_io_in_a = io_sqr_a; // @[FloatingPointDesigns.scala 65:14]
endmodule

